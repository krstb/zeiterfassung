<svg xmlns="http://www.w3.org/2000/svg" version="1.1" xmlns:xlink="http://www.w3.org/1999/xlink" width="711" height="711"><svg xmlns="http://www.w3.org/2000/svg" version="1.1" xmlns:xlink="http://www.w3.org/1999/xlink" width="711" height="711" viewBox="0 0 711 711"><image width="711" height="711" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAABkAAAAZACAYAAAAhDI6nAAABaGVYSWZNTQAqAAAACAAEAQAABAAAAAEAAAAAAQEABAAAAAEAAAAAh2kABAAAAAEAAAA+ARIABAAAAAEAAAAAAAAAAAACkoYAAgAAAQwAAABckggABAAAAAEAAAAAAAAAAHsicmVtaXhfZGF0YSI6W10sInNvdXJjZV90YWdzIjpbXSwidG90YWxfZHJhd190aW1lIjo1ODEyNDEsInRvdGFsX2RyYXdfYWN0aW9ucyI6MTgsImxheWVyc191c2VkIjoyLCJicnVzaGVzX3VzZWQiOjAsInBob3Rvc19hZGRlZCI6MCwidG90YWxfZWRpdG9yX2FjdGlvbnMiOnt9LCJ0b29sc191c2VkIjp7ImRyYXciOjF9LCJpc19zdGlja2VyIjpmYWxzZSwiZWRpdGVkX3NpbmNlX2xhc3Rfc3RpY2tlcl9zYXZlIjp0cnVlLCJjb250YWluc0ZURVN0aWNrZXIiOmZhbHNlfQBiafFxAAAAAXNSR0IArs4c6QAAAARzQklUCAgICHwIZIgAACAASURBVHic7N3NkhvXkTbgPHnOqT8UgAaaTaopybQ5Hi3IcMxiIryYjbmYW+DcDps3MRdhzXIugNpOhHcmFw5LtiUOm1ST7G4Ahfo7J/NbdBUMUrTH/ixbf+8TUYGqU9XdAESRAN7OTCIAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA+L4y3/QdAAAAAAAAAAD4C/2jPsfQf9DPAQAAgL8jBCAAAAAAAAAA8G2w+4xC9Sp/ePjw4RufWzx+/Pgrn2Pcv3//b/qhH3/88VfW7t69+0YA8uDBAyUiMuaNH4+QBAAA4FsOAQgAAAAAAAAA/D3tPns4OTl55+cQDx48ICKijz/+eHd+DDYePXq0W/vNb35jTk9Pv/I97ty58/91x548efKVtePjY/3oo4924ca9e/d0uG+7a+7fv/+V8OPhw4e7/ZOTk/3zCEoAAAC+IQhAAAAAAAAAAOCv8fZnCW8cn5yc7PbHio379+/TkydPDBHRL37xC/rNb37zxtcsFgtDRPT8+XNDRPTTn/6UXrx4YYiIzs/PDRHRZDIxq9Xqja8rimJ3fHR09Fc9iLOzM5pOp0pE9OLFCyIims1mu7Ciqiod7psSEd24cUN/+9vfEhHRe++9p0REt2/f1l/96le773l6err7+jt37ujHH3/8lWqS0YMHD/StipIRAhMAAICvCQIQAAAAAAAAgB+Wv+izgD9VrUH0Ziuqs7Oz3f69e/eIiOjZs2eGiOjmzZuGiGi5XBoiotevX5tbt27tQg2iq2CDiCjPc7Nerw0RUZZlhogoTVNTVZUhIkqSxNR1bYiImqYxRESz2YzG4+l0+pc8LMrzXImIVqvVbq3rOt0/t782mUy0bVudTqe6H5rUdb0LSJ4+fUrj/h/+8AdaLpc6PF4dng8dno83wo0xJBm9HZbshUl/TSiCAAUAAGCAAAQAAAAAAADg++td7/u/snZycvJGqLFfsfG2Z8+emf0A4+7du/Tq1avd8eHhobm8vDRERPP53BwfH9NqtTJjtcZmszF5nhsiou12axaLBW23W5OmqUmSxDRNY7z3hohovG3b1ogIF0VBXdeZrusMEVFRFERE1HWd2d9/+z4nSaJv72+32935EIKO59I01aqqKISgaZoqEZG1VoiI+r7XPM/18vKS2rbVoih0uH+7UKQsSz07O6PJZKKz2UxPT0/p8vJSh+dDX716tbsvh4eHSkT0+PFjIroKUPZDkkePHhER0dHR0W5tPyTZr7bZ864ABKEIAAD8ICEAAQAAAAAAAPjuMkR/rNa4c+eOefLkiXn27Jm5efOmWS6XZjqdmvPzczO2kKqqahdAjBUVWZaZpmlMmqa7wCFJEkP0ZqDQtq1J09R0XWf6vn8jpAghmKIoqO970/e98d6bEIJxzpkYo8myjEIIJoRgsiwja62JMe6uGX4Ej+tJklAIwYzHImKY2Vhrd/eHmd/4XENEjPf+nU+UtVaHx7PbH/V9v1uLMWqMcQw+NMaozjmNMep43LYtOec0hKDOOR0e/+54XOv7/o1r+r5X771673W73ZJzTpMk0aqqyHuvSZLoGNCMFShJkui4n6apZln2RujSNM2ueqUsS51Op/rixQuazWZaVZU65+S9997T8/NzPT091Tt37uiTJ090+HMzPg8ISAAA4HsJAQgAAAAAAADAd4chIlJVevjwoXn8+LG5e/euOT4+Nm3bcgiBJ5OJCSFwjJGdc3YymfB2u7UiwiLCqsrWWlPXNdd1zc65MVTgtm3ZWmv2w4kxeBARE2M0RMTDOR7XiYj2gwpr7bjOIrJbGwOL8evG762qu2vHY2PM7vrxWFXN/s8c7Qch++estTR8/e4DfmOM7n3dGHrszomIjudERN++NcZojJHeXnv7uuHny9vfzzkn+9cysw7hi4z7MUYVEfXei7VWjTFCRJSmqewHMuMtEYn3Xo0xwsy7bfj50Vor6/VaDg4O4suXL8U5J2mayunpqT5+/Fjv3r2rb80kQSACAADfCwhAAAAAAAAAAL79xvfv5uTkhO7cuWOOjo7Mb37zG/Phhx/yZrNhIrJVVbkYIzOz7fveEZGPMTrnnBMR1/e9DSFYZrYxRhtjtM45jjFaVeWu6+wQJnAIgekq7GAi4v21MbCIMbKI8BhOjOuqaob7Yd7eZ2YagphdqCEivBeEEBGxGT6NH6/b2+f9J2b8nvvH4/64vh+AEL0Zggyhx+7cGGiM5/Tqh+q4//b6eP27rt3fZ2Yxxqi1VlRVhvBjDD2EiGQvMBFrrTBzdM4JEQldhRxydRdFjTGSpmkMIYgxRrIsi6oanXNRVaO1NjjnQggheO9D3/chTdPQtm2YTCaBiGJZlvLFF1/IRx99pGdnZ/rkyRMd2mqhMgQAAL4XEIAAAAAAAAAA/OO8UcExLt65c2e3PwYbRESnp6e79eVyaUIIvFqtzO3bt03f9xxCYGutHQOPEIJLksTFGMfwIyEiP+x7VXV93ztVdUTkQgjOGGNV1YqIHcMOVbV0FXjY8VhEmIg4SRKb57ktisKNP3s/zIgxsjHGjCHHGIoMj3s8HgMT3ts3zLy75q1QhfbP7Yccbwcg+8b1/YCD6M0AZPgebwQi++f3g4zx/Hj9/rl3hB40hh5DhYiMt6qqQ8Ahqip938eqqmLTNCFelaOMgUg0xkRmjkQkzrlIRGKMEWNMNMaItTYMlR/RGBOMMSHLsl5EAhH1RNQ757qu63oi6r333X4goqqxbVv13svLly9lsVjoer3W169f6/HxsX700Uf6ySef0J07d5SI6OOPP97NIXnw4MH+80aEwAQAAL5lEIAAAAAAAAAA/P18JfAY53QcHx8bIqLFYmHKsjQvXrwwk8nE5Hluzs/PzXq9NlmWmaqqdgPCY4y7dlZ5njMz2xCCExFHRN4Y42kIPLquS5g5UdVERJIQQiIinogcETkR8cPmVHUXghhjWESsiNi9daarFlV2Op36g4MDf3R0lOR57pMksfthxRiA7IcVQ9DxlQBjqPzYD0bGCg6z99wZoqsP2Pe+bv/zjHd+tvF2KLIfgrwdgLy99q79/eqP4dQboch+ALK/tr/tByLWWjHGaNd1cbvd9i9fvuxev37d13Xd01XIEa21kYh2IcgQeowhSBwCkTCes9YGZu6ttb21theRTlU751wrIp21tjPGtETUG2PGQCQ0TSMiEplZyrKMm81GnHMynU61aRqt61qrqtJ3hSNnZ2d6//59JSJ6+PAhoZUWAAB8myAAAQAAAAAAAPj67YaT7wceY9iR57nZbDZ8fn5u+r7n6XTKfd9znuccQuCmaczYXkpEOEkSjjE6EeGu66yIOGa21lpX17UnIq+qybgRkReRlIhSIkpUNYkxJqq6qwQZQxMRcWMIMoYeNIQde2u7NljXr1/PPvzww/yf/umfisVikeZ5vps6vle9Qe8INGjv+I3Q4+1z7/h6etd1X5d3BSJvn3vHNe9sq/Wu69+uINlf22634fz8vP3000+3T58+rV+9etXSVQVIZOY3QhAago8xEGHmMAYlw1qw1nbM3BtjemNMR0SttbYlolZVO2ZumLlj5o6IehHpmDkwcxhaaAVrbcjzPLZtK6oaQwhqrZXZbBb7vtc0TaVtW83zXOq61rIsZbPZ/LlB6whCAADgG4EABAAAAAAAAODrY05OTsyDBw/o448/Nufn57xYLExVVdx1Hed5/kbgYYyxIQQ2xthxIyI7Bh3j2hB+7La9ECPx3id5nqdZlmXW2pSIEiLyfd8nqpqObbBExIcQxoqPN76fqtphDsgu7BjCl6+svffee+n7779f3L59u1wul2lRFH7/CfgT4cQ7P3/4c0HG/xVyfJ0hyJ8LQL6Oa95e3z/ebrf9+fl597vf/W7z+eefb8cAZGhvFYloDEF2bbHoamB6fCv8iGOQwcz9XiVIO4QdHTN3qtqoats0TdN1XdP3fUtE/RiIeO97IurHGSKqGokoElFU1aiqcTKZxKZpxDkni8Uibrdbuby8lCzL5E+FIXuVIQhDAADgHwYBCAAAAAAAAMBf7p3vo09OTt6Y57EffFy7do3ruubz83NrrbVFUTAR7cKOvu9djNFZa12M0TGzezv0oKsAI4kxeiLyIYSx0iMtiiKbzWbFcrkskiTJjDHpEHD4EEJCQ7urGKOLMb5R6TF8f6uqvBeAmLHllary3r4RET48PEyPj4+zDz/8sDw4OEj2K0Dgr7fdbsPl5WX39OnT6tmzZ/XFxUU7tMoSZhb648wPGdfHmR/DEPUxEJG9EGTXDssYMwYhnTGmV9Wm67pmtVpVq9Vqu16vaxqqQ7z3Y3VIS8P8EGttoKFl1hiIeO9DkiRhqEqJMcZQ17WoakySRM7Pz+Wjjz6Suq51f8g6EdEYhhDt5oaMEIwAAMDXDgEIAAAAAAAAwLv9X5UM5v79+3R2dmbu3btHz549M//6r/9KbdvydDo11lp7cXFhp9MpM7M1xti+711RFNZaOwYUbmhL5YwxyVitYYzZhR7jFmNMiSiNMaYikopIysz5YrGY3LhxY/bBBx/MyrIsvPf+rRkeuyHmw5oZg43hHI9tqvYHl781r2N3m+e5K8vSLxaLJMsy5723f///FN9ffd/Huq7j5eVlt1qt+rZtw/7cELoKQN6eJ/LGcHVV3Z8vsh+WjJUhuyqRvu/b7XZbP3/+/OL58+fr169fr1W1NsY0zNxYa2vnXK2qnTGmHVpqtUOQ0nVdF4b2Wr1zLjBzH2MMIYSQpmmo61pEJHrv5fLyUpxzkiSJ7M8OGStDxoHqJycnRO8OQBCKAADA3wQBCAAAAAAAAPyQ7WZ1EBE9fvzY3L171zx79szcvHnTLJdLQ0T0+vVrc3l5aebzuSEi2mw2ZrvdmrIsTVEU5uLigrMsM1mWGSLiyWTCVVU555wdJUniRMQZY7xzzo0Dy0UkGfZTY0xijPEispvnoaoJM6fOudx7n3vvM1XNiShV1WKxWJQ3b96cvf/++4vpdJp77z3tBRbj/n6YQfSn53Xst5Z61xwO5xx774333lprDb89bRz+KjFGFRHpuk5CCBJj3E1r3x+4vr/2p+aNDIPY96/Z3RKRMrN0XddVVVWfnp6ev3jx4vL169crY0xNRI2qbvu+34YQqhBCLSItEbXj3BBjTBtC6EWko6FCRFV7Ve1DCIGZQ9d1IcYYkySJdV1LkiRxu90KEclsNpO2bdUYI0VRaF3XWte1bjYbLctSZ7OZLhYL/cMf/kDL5fIrgcn9+/cVg9YBAOCvgQAEAAAAAAAAfmiMqtLDhw/NGHiMA8qfPHnCx8fHu1kdIQSOMXLTNGN1BHddZ2hoDxVCMKrKbdtylmVMRBxCsDFGa4xx1lpLRG7crLXeWuuY2atqYozxzOxDCIkxJnXOeVVNRCQhosQYkxBR4r3P8jwv5vN5MZlMiiRJ8mHIeT6fzyfXrl2bHR8fz8uyzIYABOCduq7rt9ttc3Z2dv7y5cvVxcXFxhjTEFHT9/12s9lsLi4u1k3TbEMItTGmE5GGmVtV7WKM4/D0XfgRY+yMMX0IIRBREJE4tOYKNMwtCSFEIpLJZDIOc5eiKMQYIyEEzbJsHLCu1lqx1or3XsaWWovFQsuylOvXr8t6vX6jpdYwaJ0IYQgAALwFAQgAAAAAAAD8kJiTkxMzzulo25ZDCHzt2jVmZts0jRvbVYUQnDHGbrfb/TU7BhwxxnF+x67dFF3N27AxRjcOHCciN5zzROTG9lZ0FYrs3ybj8RCQeLpqh+XzPE+Pjo6KW7duTW/evDmZTCYZMydE5NI0TSeTSVaWZZ6mqR9CF4B3CiHEvu/7qqq2VVU1bdu2Qxurrqqq+tmzZ+vf//73l69evarqum6JqBORbgg7OroKOHpmDjHGYIwZK0ECEYWh1dbulpmjqgbvfdybTRLzPA/W2qiq4yD34L2PzrmoqtE5F6y1IUmSkKZpIKJdG68syyRJknh2dibjsHUiEgQhAADwNvdN3wEAAAAAAACAr9HYsomIaFflQUR0dnZmPvroI/Pq1St++vQpxxg5TVN748YNOwwd95PJxImI77ouERFvrXX+qteTa5rGj8PEicjFGL2qji2txs0ZY8aB434cYj5uxhi7t+9ExKmq3dt3dBWSWLoKThwROedckqZpMZvNpovFopzP59kwe4OZ2XrvrffeMTN+0RH+LGutISJXlmWRpmkaY4zGGIkxBu99vV6vJ0mSZNba7dD2qjfGBCIKqtobY6KqhjHk2N8fb40x0Vr7RhDivQ/jYPYYY6+qXQghWGv7GGOw1vZ93++OiagzxvQxxq6u636cNZIkSWDmsN1uQ5qmMc9zmc1m4pwbAxB5/Pix3r17V4mI3jFwHeEIAMAPCF4YAQAAAAAAwHfZGzM8iIiPj48NEdFisTDPnz83IQSeTCbm9PSUl8slxxi5rmu7WCxskiTOOef6vk/GigtmTlQ17fs+HVpR+WEA+S4YiTEmIQQfY/TMnKRpmh0cHKSTySRLksSrqhvOj4GHVVUbYxwHk9uhpdYbg8qHSpHdvjGGVdVlWeauX7+e/eQnPyk/+OCD4uDgIHHO8f5zsPcBL97rw5+jRH8MCcfjEIJcXl62//u//1v99re/Xb169app27Y3xkQiiqoax3CDrlpYRWvtbn8IOmSo5tjtM/NYzRGZOfR939V13VxeXtZt27aq2jFzb63tnHOdqvbM3FlrW+99Ow5iV9VuqEDpxyHsSZKEzWYTRSTGq0ns0VorzjlZLBZaVZWOw9efPXumN2/e1MePH+vHH38s+48dAAC+v/CiCAAAAAAAAL6r3mhntVgsTFVV3HUdhxB4Pp9z3/dcVZUVEbbWWma2MUYnIm6s1vDe+67rUmZOQggpXQ0XT4cZG6mqJjHGNMaYDMPJfQghjTH6q1nPSbpYLIoPP/xwcv369WJoT2VFZAw5WER43B8GjbOIMF3NI9mtqer+2m7fWmvLsvRHR0fpYrFI8jx3GD4OXycRkbquw8XFRfvy5cu6qqo+xhjpKiQQY4wMt2qMkWG4ujCzMLPQMHCdmWU8P4QhundNqKqqOTs7q54+fbparVZ113Wttba31rbW2s4Y0zFza4xpnXMNEbXOuVZEWmbuVLWz1nbjIHZVjTHGoKq9cy6ISMzzPNZ1LWVZRu+9rNdref36tVhr5YMPPojn5+e6WCzkyZMnSkQ0VI4gDAEA+B5CAAIAAAAAAADfNWb47XXz6NEjPjs7YyKyTdO8c45HCGHXgmqo9vBE5L33XkQSZk6MMRkRZc65jJnTGGM2BCCJiKQikoYQUlX1McZkqABJYoxJlmXp0dHR5Pbt27MPPvignM1mmbV2DD+MMYaGgMOoqtl7DLvjcZ+ZaX9tvM5cJTWc57lNksQ659jslXwA/K1UVUMI0nVdrOs6hBBEr/7wKQ3hho7/412t0RCGjOfeON4/P+6LSFitVs2LFy9Wn3766cX5+XnVNE3rnOuYuXPOtWP1hzGmsda2zNyMgYgxpo0xdiLS9n3f9n3fOed6Iur7vu+9932apmNLrRBCCKoavfdBVWPTNOHHP/5xGOeHHB0dySeffEJEJA8ePNjdVwAA+P7AiyUAAAAAAAD4Lti1unr8+LG5e/euISK+desWW2ttlmWurmvnvXdN0yRE5FXVj4EFXbWxGis4EmNMEmPcVXnkeZ6XZZlPJpMiSZLUWpuFEHYVHzHGdBhqngwVJMlQAeLGCpAf/ehH0+Pj43I6nabOOd4LO4hoF2hcPZi3sou3r317fbjeWGvJXNk9JwBfE1VVUlUVkXGf/lQo8Pb62FLrz10fY5TNZtO8ePFi/cUXX1xcXl7Wfd+3zBzGFlhDFUhvrW3HQGQIRboYY9v3fbPZbOr1el1vt9t2mFPSqWrnnGuttd1eO62OmXtm7ofKkd4512dZ1r98+TK+fPlSnHOSpqm8NUgdQQgAwPcEhqADAAAAAADAt83bH+ybk5MTGoaZm/v373NVVbuWVkmSOCJKiChp2zZ1zqVElA1VG9mwnxFRSkQZEWUxxizGmKlqpqqZc24ynU4nx8fH5WQyybz3qYg4IrIhBKeqTkTG9lnjPA8nIuycc3mep8vlMs/zPPXee7Sngu8gY4whY4z5e/3xNcZIlmW8WCyYiNzR0VEXYwzMHIcB6dFaG4wxYQhF+nGIOjOHruvaqqoaVV1XVbURkXpojdUyc0NEjTGmds41xpjd5r1vrLVNCKFxzrV937eqGiaTSQghRCKS5XIZf/3rX5t79+7pvXv3hOgrA9QRigAAfAfht0UAAAAAAADgm7ZrC3VyckJ37twxT5482X+/yq9evTKHh4eGiPjo6Iidc3axWNjLy0u/XC593/dp0zRZjDFn5twYk4cQClXNRWTCzAURjcd5jDEXkVxEMhHJr127Vh4fH5c/+tGPZvP5PMuyLKG35nOMMztEhI0xZq/F1ViFMg5VR3sqgHcY22z1fR/atu1jjKKqMswN2c0WGW53m6qqtVbquu5Wq1X9xRdfXJ6enq5ev35dDUPSG2ttba2tvfdba+1WVbdEVKnq1jlXWWu3fd/XRFQTUT0OVV+v17sB6m3bRmut/O53v5PDw0M9Pj7Wjz76SD/55BO6c+eO3r9/Xx8+fDjODCFCKAIA8K2HF2QAAAAAAADwjzTOt6CHDx++McD8yZMnfHx8zCEEjjFymqYmxrgbIL4/yFxEnDHGE5EnotQ5lxpjshhjEWMsRKQwxhTW2iLLsrIoijJN09JaWxBR1vd9Pg46jzFm8/l8cnR0NPnggw/K6XSa5nnuh/u5m8cxzvLYXx8f0/Bb8+Pt7nECwBtUREiviIgQDSHC/qyQ8dq31+u67quqak5PT1dnZ2fri4uL7dDyqmXmxjnXDOFH1bbtpqqqVdd1VYyxIqItEVVD1Ui9N1MkhBACM4ftdhtDCDFN0zgObl8sFrLZbMQ5J9evX491Xevz58/l3/7t32S9Xo/VIooqEQCAbye8IAMAAAAAAIB/FHNycmLGCo87d+680cpqHF7e970LIThmtsxsY4xuPKeqzhjjQwheVcd5HqmqZsycxRhzVS1UNSeiPE3T4uDgYHr9+vX5crmcZllWGGPSYb6HjzF6EfFFUWTz+TxbLpd5URR+aKsFAN8ifd+Huq678/Pz7Wq1qrfbbTu0yQrDzJCOiNqu66qLi4vV6enpxWazWXddt1XVLTNvhwCkIaKWiFpV7b33HRH1McbgnOtDCME5F5k5FEURxiHqzNwTUVTVWJZlODo6Ck+fPo1HR0dy7949QXUIAMC3DwIQAAAAAAAA+LtTVfPw4UNDRHznzh0uy9LEGK2I2IuLi0REPDMnfd8nw2Dy3fDyrusSY4yPMe5CDxHxIpKKSKqquxkfY0srVc1VNU3TtHjvvfemP/3pTw/ef//9eVmWhXNunOPBw2attTZJEptlmXPOWWstZngAfMuIiAytqkLXdSHGGIlIjDHCzNEYE1W1X6/X29PT04tPP/309atXr9Z1XW+NMS0R1czcGGMaVW2ZuTXGdMaYbtwnot4Y01lre2buvPe9MaZ1znV5nrdE1A2hS5ckSe+9727fvh0uLy9lvV7rf/7nf+rdu3f1wYMH+qcGwgMAwD8OAhAAAAAAAAD4uhjaG1h+9+5dQ0R0fHxs2rblEAJfu3aNLy4urHPOZlnm8jz3fd+nMca07/sshJAZYzIRyVQ1VdUkxjgGHYm1NsvzPC/LMvPej0PMkxBCKiLJsKUxxkREkiRJ0sPDw/LWrVuz9957bzqdTjPnnH2rldWuhdXYxgozPAC+ffSPvbN2LbSGkEGH2SEaY4zr9br58ssvV59//vnFxcVF1fd9MwYdQ7jRGWN6a23HzB0RtW3btnVdb9u2bdq2bY0x3TA8fZwx0jBzba1tDcqx0QAAIABJREFUiajJsqwRkdY519R13atqvLy8FOecJEkik8lEzs/P9fT0VImIHj9+rHfv3lWiq+HqaJkFAPCPgRd0AAAAAAAA8LcyJycn5vHjx2axWPDNmzfNcrk0IQSeTCYmhMDOOVtVlR2qKywReWOM996nY+gxVG3kMcZi2M9UdQxF0hBCWhRFcXh4WB4dHZVFUeRJkqQhBD9UhLihrZUb9p211k+n0/zGjRvFYrEoiqJIUN0B8P0VY5SxTdbLly/X2+22CSH0xpjAzGFolzXe9swc+r5vq6pqzs7OVpeXl9u6rrfM3DJzzcwNEdVJkmyttVsiaqy1taqOs0S2ItKNbbJUNVZVJbPZbBeIVFWlzjl5/fq1Hh8f6+npqY6ByNAyC0EIAMDfCQIQAAAAAAAA+P82VlA8fPiQiYhv3brFL1++tMvlkkMI3Pe9G2d8hBDcOLw8xphYa5Mx+BCRgpnzGONEVSeqWgytrDIRyceKkMViUd68eXP+4x//+GA+nxd5nmeqyvstrcaB6UTExhhOksRlWebzPPfOOcvMeC8M8D0lIjq0yerruu5CCIGIIl1ViQgNLbOGtllijJG6rtvLy8vt73//+9dffvnl+vz8fGOtbYwxtbW2ZuaKmbfOuUpVa2vtNsa4ZebKGLMNIbTOuc5aG0IIQVWjcy6oahSRGGOMzjnx3kuWZfL8+XNJ01QWi4U8efJET05O5Bt+2gAAvrcw1A0AAAAAAAD+amPw8ejRIz47O+M7d+7Y9Xrt6rp2h4eHru9757133nvfNI0XEd91XWKtTYbZHqmIZHmeF3meTyaTScHMhYgUMcYihLALPWKM2dDWKp3NZpPFYjGbTqcHs9ksz/M8He+LqhpjDKmqGTciMtZaY63lqxwGxR8A32fMTM45HirMrKoK/bHCYpzLoUS0a5/lnOtEZHtwcOBjjBPnXMXMrXOuds41zFw752pr7dZaWxtj6hDCtm3bzXa7XccY667rWiLqrbUdEfWq2llrd0PVvfchTdNQFEX46U9/Gl++fBmrqoq/+MUvgqru3zcAAPga4bdeAAAAAAAA4K9ycnLCd+7cMbdv3+b1em3Pzs5c3/c+xuiZeZzHkYYQkhBCRkRpjDEbZnlkY1WH976Yz+fle++9Nz04OCizLCtUNRuuHed5JDHGJMboRcRPJpNsPp+XR0dHZVmWWZZl/pt+PgDgu61pmr6qqubLL79cr1arbdM0NTP31tpumBPSWmtb51xrrW2NMU3TNNvLy8vV8+fPL9frddX3fW2MaZm5YebGe98Ox61zrvPed2madm3bdpPJpGvbtt9ut32SJP3t27fDf//3fysRydASiwhtsQAAvhaoAAEAAAAAAIC/lDk5OTF37twxRGQ/++wz23WdL4rCxxhTIspUNSOi3BhTWGvzGONERApVLYhobHFViMjEWlt672fT6XR+/fr1aVmWhbXWi4hTVSsidmhtNd6yc84lSZJMJpPEOYdyDgD4mznnuCiK5Pr16+XBwUEaQpgOLbIiMwdmjsaYyMzBWhtijH1VVdsY46X3/hURrUWkGmaDbIloG0KonXM1EW1jjI1zrh7XQggNM7dJkjRlWdJnn31Gy+VS0jQ19+/fl2E2yHj3EIQAAPwNUAECAAAAAAAA+wwR0TjU/O7du+b4+Nj8+te/5sPDQzOZTOxyueS2bZ0xxotISkQpM2cikhtjCiIqVHVCREXXdVNmnjjnyjRNJ865kogmMcYiSZLJcrmcffjhh7MbN26Uk8kkH1rW8H5bq/F2aHHFzGydczzA+1oA+JuIiMowrENERFVlbI+1dyvGGDXGSAghbrfb+ssvv1w9ffr09cXFxSaEUFlrG1XdhBCqrus2McZKVStmrq2126GVVqWqtarWzLxt27ZxzrWqGpumCSGEeHR0FMc5Iaenp0pE8uDBAzVm99cdQhEAgL8QXigCAAAAAADAaFfhcX5+zqenp/b4+JgvLi5skiTWe29DCI6ZvTHGt22bWmszIsqJKBeRwlo7McYU4zDzEMI0SZKyKIrpYrGYFkUxS5JkEkLInHPFdDqd3Lhxo7x27VpRFEVqrUVVBwB8q4lI3G633atXrzZnZ2eXVVVVQ5VH03Xdpmma9fn5+appmk3XdRtjTM3M22GriGhrra2IaGuM2RJRo6odEfXGmJ6ZexGJIhKHge7xZz/7WTw7O9NhaPpujgkAAPx5CEAAAAAAAACAiIjv379vFosF37x5096+fdvGGL2qelX1zJz0fZ+oatp1XRpjzEIIOTMXIYRCVYuxtdWwn4tIISLFbDYrl8vl7Cc/+cn82rVrs7IsCxHxROS898lkMknyPPfee4eKDgD4tlNV6fs+1nXdbbfbNsbYqWqw1obNZlO9fPly9cUXX5y/evVqU1XVZpgFMg5Sr4ioNsZUxpjKe18557ZE1IzbMDekFZHOWtsfHBx0L1++jNeuXQtffPGFLBYLGYIQ+WafCQCAbz+8sAQAAAAAAPhh2b0P3G9zRUR8eXlp5/O5JSJXlqWbTCapqqbe+7Rt29wYk6lq3nVdEWPMVbVwzpXOuUmSJKW1NieiIsaYi0gWQshEJJtOp8VyuZz+5Cc/md+4caMsyzJXVR7aWbG1dmxpZcxejxcAgG8jVVUR0ThQVSEiUVXdbDbbly9frj///POL169fb7bb7ZaIeufcGGxsVbU2xmy7rqv6vl+LyJaItt77ipkra20tInWapk0Ioe37vs3zvGvbNmy329C2bfzggw/i+fm5jmHIgwcPlIhoaNkFAAADDEEHAAAAAAD44TD3799nIqIx9Lh79y4TERMRz+dz17atT9PU932frFar3DmXtW1bGGOKYb7HRERKVZ2IyISZZ3mel7PZbJqmaW6tzUMIaYwxEZEkxphMJpPs4OCgmM1m07IsJ2VZpt/kkwAA8LcwxhhrrRla9vn9c6rq27Z1y+XSGmOKoiiaYXh6Z63thsqOuu/7er1eb2KMq77vN8y8adu2staumLli5qqu6y0z10RUX15etiGETlX7LMvCer0Oq9VKqqqS5XIpjx49imdnZ6qq+7NLAAB+8BCAAAAAAAAA/ACcnJzwo0ePdoHH8fExn56euqZpbJZlloicqibWWk9Eadu2WZIk+RByFKpaGmNKIprGGMsY41REyul0Ojs4OJh98MEHs7Is8zRNsxijExGrqlZEnPfepWmazGazzHtvv9lnAgDg78d7b6fTaUZEtFgs8hBCz8zCzNFaG4wxoeu6drvd1s+ePVvXdX3Zdd3aGLNm5rWITJl5bYxZE9GGiLYiUolIQ0QtEbVd1/XW2r4sy1jXdSCisNlsQlVV8qtf/Sp+9tlncnJyglkhAACEFlgAAAAAAADfa6pqHj58aOiqysMdHR25ruuctdbXde37vvchBB9jTGOMqaqmxpgsSZI8TdNJlmXToihKZp4SUSkiYwBSxhgnh4eHs+Pj4+mtW7dm8/k8y/M8ERFWVUNERkTYGMPOOfbeW+ccY9A5AHxfxRglxhhDCDGEICKixhhlZqGhMqNpmm69XjdPnz5dP3/+fHVxcbFm5g0zb5xzl8P+WlXXbdtWdV2vt9ttTUQ1MzfD1g1tsfqiKNrr1693IYTQ932oqir87Gc/i5999pncv39fUA0CAD9k+M0bAAAAAACA7yFVNcYYPjs747OzM75165abzWY+y7K07/u8bduCmScxxikRTUVkpqoLIlqIyIKZl1mWHS0WixuLxeLGwcHBjclkclQUxVFRFIdFUSyLolgeHh4uDg8PF0dHRwfT6XQ6mUwmaZpmWZalWZaleZ4nWZb5JEncOOfjm35uAAD+XpjZWGvtUPnmsyxLsixL0itZkiQZM6dElHRd50Ukcc6lZVlmZVlm0+k0n81meVmWkyzLCiLKq6rKuq7L+r7PjDGZiGTOucRam6Rp6qy1VkQ4hMAiYpiZ+r43IQT6r//6L3Pv3j169OjRN/3UAAB8I9ACCwAAAAAA4PvFXLWAJ3N8fGyfP3/Os9mMvfd+vV5nqpozc2GMKUSkEJGJqk5omO0hIpO+73Pn3CRN09n169cXN2/enJdlWTJzFmNMxk1EkjRN06Io0qIovHMOlR0AAP8H55zJ89wfHR3leZ5z13WptbZk5s573xhjOiJqNptN9eLFi9X5+fl5jHEjIhsR2SZJshGRrYhUIYSKiDYhhI33vk6SZOucs6vVqosxmp///Ofhf/7nf+jk5EROTk7Gu4CKEAD4wcBv3gAAAAAAAHz3GboacG7G4ea3bt3ily9f2jRN7eHhod1sNlnbtgURlXstrKYiUsYYZ8w8U9WZiJQhhDxN08mNGzfm//zP/7z48MMP5/P5vLDW+mGuhyUiFhHLzDZJEk6SxFprmZkRggAA/BkiojFG6bou9n0fRSQyczTGiDEmMnOMMfar1ap+9uzZ5aeffnr+6tWrdQihStO0stauiWijqmtjzMpae+m9X1lrN977ipmrrusaZm6cc/0f/vCHUFVVJCIhInn8+LHevXsXM0IA4AcBAQgAAAAAAMB3lzk5ORnne/BsNrOr1coeHx/bvu9d3/dJ27Y+TVPHzEUIoTTGzEII0xDCTESmzrmZ934+mUwWaZoeMHPZdV2WJEm+XC6nt27dmr///vvT6XSaOefeaKM8zPkgYwwZs3t7ifeZAAB/nhIRDdV6pKr09pyOGGNcr9fNixcvNr///e9X6/V6E2Pcpmlai8i667rVdru96Pv+UkQuvPeX3vuVc24cqL5V1bqu685a2zJz3zRNCCHEoijCZDKRo6MjOTs7U8wJAYDvM7wwBQAAAAAA+O75SvAxn8+dqvq2bRPnXNI0TRpjzEQkE5GMiCYxxulQ5TGNMU5jjNOiKGaLxWJ+8+bN5cHBwUGe55MYoyeiZDKZpMvlMp/P53mWZR7VHQAA/xgiIk3T9KvVqj0/P9+2bdsSUeec65um2axWq8vT09Pzy8vLy7quL5xzK+/9OkmSFRGtmbmy1laqWltr6yzLmiRJWmNMt1wuO2NMOD8/j9bamOd5/OSTTwQVIQDwfYQZIAAAAAAAAN8hJycn/PjxY/Ps2TO+efOmvX37tq3r2hljEmNMZq3NYoy5MaYwxpTGmCLGODHGlMw8M8bMVLW01pYhhDLP82lZlvNr164tb9y4MZ/NZoWIMBGxtdZlWeaSJLFmr8QDAAD+vowxxnvvZrMZpWlqRaQgIjHGyGazqay1k9VqlTVNM+n7fuK9nznnNsy8VtVVjHGjqushBNnEGLdEtGXmZr1e133f99baLs/znq5mRsVf/vKXgmoQAPi+wQtYAAAAAACAb79dxcfx8bFp25Y///xz96Mf/cgWReFijCkzZ23bFsaYIoRQxhhLEZmFEEoRmSZJMk3TdF4Uxdw5NyGiSQghL8tycnBwML1169b8+vXr0+l0mqnqmHcYZjYDIryHBAD4R1FVJVVVEdlVZhhjdL1e169evaq++OKLy4uLi01d12vv/dYYU6nqpq7ry7ZtVyKyZua1c26VZdmaiKokSSprbdU0TcvMDRF1i8Wia5qmt9bGL774Qk5PT5WI5MGDB4owBAC+6/DiFQAAAAAA4NvpK4PNZ7OZjTFyjNGVZemMMb7v+8Q5lw2VHtMx+IgxzkXkIMY4izHOZ7PZ7PDw8ODGjRvzyWRSeO9zEfHe+zTLsvzw8LCYzWZZnuf+m37gAADwpzVN063X6/b8/Hxb13UTQmi9923f93Vd19WXX355sVqtLtfr9Tgg/SJN0xUzr7z3677vN+OMkCRJ6hhj23Vd2zRNyPM8ZFkmRBTHGSFPnjzBwHQA+M5CCywAAAAAAIBvH3P//n0eg49bt27xdrt1zjnb9/0u+BCRJMaYEVEeYyyH9lZzETlg5gNjzMIYM2fmgzRN57PZ7OD69euzxWKR53meqiobY5xzzqZp6r33mPEBAPAt55yzZVmm3nuOMeaqGpk51nXdrlarbVVVk+12WzLz1Fo7McYUqlqEEPIYY6aqKTOnMcZ0+Lekds65JEk6Ve2JKMzn80BE8e7du3J0dCS//OUv9T/+4z+EEIIAwHeM/abvAAAAAAAAAOyYk5MTJiL785//3M5mMzebzXwIIe37Pk/TNG+aZjJWeYjIXEQWXdct27Y9DCFc895fK4ri+sHBwY3ZbHa9LMtrRVEcLpfL5dHR0cGNGzfm8/m8nM1mRZZlaZZlyRB+WGstY9YHAMC3mzHGMDN7712apj5N0yRN05SZvTHGN01jr0aI+GQ2myVlWSZZlqVElHRd59u29X3fpyKShhASY0wSY0yMMd4Y47Mss33fWxHhV69ecd/3HEKgu3fvmnv37tGjR4++6acAAOAvhgAEAAAAAADgm2eIiO/fv8//8i//Yq9du+aIyGdZlnjvM1UtmLlU1WnbtnMROQghHPZ9fxhCuBZCOOq67khVr6dpeuPw8PDGjRs33rt27dr15XJ5OJ/P58vlcrpcLsuDg4N8MpkkSZJ4e4WttTzO+vimnwgAAPjzhgDEjH9/D3+XWyLicUvT1JdlmS6Xy6wsyzxJkrzrunS73aZVVWUhhCKEkKtqoaoZEaXW2tR7n9DVvz9WVS0RMTOboijIWmuKoqA8z+nJkyf49wIAvhPQAgsAAAAAAOCbZ+7fv2/+/d//nauqcnmeu8PDQx9jTLuuy9I0LVS17Pu+9N5P2radhhCmqjoVkWnbttMY4yTGWDLzfDKZHBwfHy8PDg5K730qIm7g8zx3zjm0ugIA+J5xznFRFP7o6GiyWCzSEEKw1oau65r1er3dbDYHqnrRNM3KGLOx1lZEtGHmtYisVHVNRGtm3sQYV865iv4fe/fSI7eZ3Q38PDc+vLNI1q1b0ivbMCYTKUAGCDBbezHLySaADOQLZJEPkK0rX0faZj/yIgiQLCZAYA0QBDMe+CJZfa0ri+RzeRfd1dNqt2TP+KLb/wcUqppVxSJbra5q/nnOIdpIKbn3njnn+rIs2a9+9StDRO7BgwdEaIkFAK84pLUAAAAAAAA/HUZENJvNGBHxvb091rYtPz4+FlVVSSml2M33MMaERBRJKSPGWGqMya21mTEm9d7nQRAUQRAUSqmCiNLzPvBxWZbprVu3snfeeScviiLWWsvz1+XnZwyznZf4fQAAgB+YP2et9d57T0SOiPx2u+1Xq9X2888/Xz558mR5fHy84pw3SqmNc25trV10XXfqvV8wxhZa64UQYsEYW2qtl865jXNuY4xpnXOdEKLfbrcmyzLz5MkTp7V2jx8/9h9//LEjIn/+9oJgBABeCfjACwAAAAAA8NNgu+CDiHie50JrLbquk0IIZYwJoihSbdtqa23onIs55zERJefVHrlzLjPGZEqpLEmScjgcDoqiKKSUqfdeO+d0kiThaDSKxuNxkmVZEAQBWh8DALzF+r436/W6f/r0aXNyctKs1+uGMdYJIbZd123W6/X8+Pj4pGmahXNuobVecM7ndFYNshBCrIUQK+99Q0RbY0wrpWyFEL2Usiciu7uMRiP3ySefuNls5l7qTgMAnMMHYQAAAAAAgB8fu3fvHjfGiNu3b4vBYCCDIAi01qFSKhZCJM65zHufW2sHfd+XzrmL+R7OuaExZmSMGTrnaiHEMM/z0f7+/uTmzZujvb29ajQa5aPRKKnrOh4MBjpJEqWUwlBzAAAgIQRTSok0TVVZlno4HEaDwSCO4zi01gar1Uo2TRMYY3YhvHbOhd57bYwJGWPaWquFEAFjLOCcy7PVCpGmKffesyzLqOs6ev/99+ndd9+lhw8fogoEAF46fBAGAAAAAAD48Xyj6qMoCtm2rRRChJzz0Hsf930fO+eSrutiKWUqpczCMBwEQZByztO+7xNjTOqci621kZQyKcuyuH37drG3t5elaRoKISQRXQzGlVJisDkAAJD33jvnvLXWWWudc84zxry11qzX6+3XX3+9+vzzz+eLxWJljFkrpTZKqRXnfC2lXBHR0lq72G63S+fc0jm3VEothRAbKeVGSrn13rfW2naz2fRBEPQnJyemLEv36NEjP5vNPKElFgC8JBiCDgAAAAAA8MNjs9mMffrpp+yrr77i+/v7YjQaya7rJGNMMcYCIUTUtm3KGMu891nf97n3PpVSDrIsG4zH4zqO40JKmfZ9HzrnQmutNsZoIUSYpmlc13WSZVmcJEkghMBgcwAA+AbGGBNCsKvvE9ZaxxiTXdeJrutknuexc24rhOiUUo0QYiuEaIwxq7ZtT8/bZJ1Ya0+ttaec82Xf9yvn3IZzvjbGSM55u16veRRFPE1Ts7e35+7fv+8ePXrkP/74Y88YQxACAD8ptMACAAAAAAD4AXnvd1UXfDweC+ecLMtSaa1VFEWac66dcxHnPHPOFc650jlXOeeG1tpRkiSTwWCwf+vWrduj0ejGaDTaq6qqLsuyrOu6qKoqr+s6LcsyzrIsjKJICSHQ6goAAP4STErJ4ziWeZ7rsiyjuq6TqqrSsiyLwWBQRlGUnYf2wXa7DbbbreSccyLi3ntORNwYc/EepLUm7z1JKZlSitI0Zc459vvf/57u3r3LHj58+PL2FgDeOviADAAAAAAA8P2x2WzG7ty5w05OTngQBOLw8FBYa6WUUmmtAyLSRKQ556ExJk6SJA+CYKC1rhljA+dc2bZtkaZpWdd1dfv27Wme50UURbH3nnvvGZ0dbGJExDnnXErJhRBodQUAAH8Jb6311lpnjHHee0dEnnPuGGOOiDxjzDVNs1kulydPnjw5nM/nR+v1+jgIgmMhxCkRnTZNMz+/rLz3ayFEwznfeO+7KIq6vu9NmqaGc27/8Ic/WK21e/z4sUVrLAD4KaAFFgAAAAAAwPdzMefjyZMnYjAYyDAMpfc+aNs28N5r51xkjImdc/H5HI8kiqIyiqKqqqqhlLIkokHXdWkURUWe50WSJMM4jtMwDKOXvYMAAPBGumiNFQTB8x/EmDbGyDzPpRAiPH9vyolo3vf93Dl3vFqtTrqumxPRyjm3FkKshRCNc25LRK0xpkuSpK2qyqzXa0NE7P79+/ajjz7ahSAIQgDgR4EzhAAAAAAAAP4yjIjo/v37/NGjR+LOnTui6zrFOQ+cc+Fms4mJKLbWJsaY1Fqbd12XOecyY0y2t7dX37x5c3jr1q1xkiQDpVRqrQ2EEFpKGaZpGiulAimlesn7CQAAbzFrbd91Xds0zdYYs/Xeb6WU277v16vVavH5558ffvnll0eHh4cnQoillHIphFhorVdRFC0ZY2sp5cZ7v0mSpFksFu12u21PT0/N8fGxnc1mjhCCAMCPBAEIAAAAAADAd3dR7bG3t8fatuVaa9G2reScqyiKdNu2YRAEcdd1KRGlbdvmxpjCez8QQuRCiEIIke/t7dX7+/v1rVu3RmmaZlrryDknOOeCMSaklJJzLs77rAMAALwU7ox1zhnnnCUiS0S27/tmsVisv/zyy6PHjx8fHh4enlprF9baBRHNpZTzMAwXRLRUSi2FEEvn3MZau7HWNtbabrPZmLZt7R/+8AdX17X99NNP/d27d/15eywihCIA8D0hAAEAAAAAAPh2F8EHEfE8z8VisRB7e3ui73uplAq6rgs556H3PnLOZc65jDGWt21beO8H3vtKKTVI07TI87yYTCbVeDwup9NplaZprLXWL3snAQAAvqu2bbv1er15+vTp6ZMnT04ODw/nm81mvt1uF23bnggh5lLKuVJqzjlfcM7nzrmVEGJljNkYYxpjTKeUMmEYGuec/f3vf2+JyO0umBMCAN+XeNkbAAAAAAAA8Ipj9+7d43/7t38rOOcqz3OllNJKqcg5FzVNk3Zdl1tri67rBn3fV13XDY0xddu2Q2tt3fd97b0fJklSD4fD4c2bN4eTyaSqqipLkiRSSilUegAAwGvGM8YY51wopWQQBMoYo5qmkZvNRlprFREpa23Q931gjFHe+8B7r9q2DRhjSmutGGNKCCG99yLPcxYEARuNRvS73/2O/v7v/94/fPgQAQgA/MUwBB0AAAAAAOB6jM4qP3hVVWKxWEgppeKcB23bhowxzRgLvfcJYyzlnCdJkuRKqYwxljvn0q7rMu992vd9LoTIB4NBUdd1MZ1Oi7Is4ziO9XmrK4QfAADwWjkfnq6KouBSSqmU0m3bBk3T6L7vQyllIoTIpJRLzvmKc74QQiyccwvG2NJau/Ter4UQDRE1YRg2XddtOedd13Xtr371q+7k5IS890RnYQuCEAD4s6EFFgAAAAAAwLMYEdFsNmMPHz7k//AP/yCEEIoxptq2DcMw1OeDzWPvfeKcS4loEEVRUVXVIIqiQilV9H2fWGtjY0xsjEmIKB0MBul0Ok1v3bqV5XmugyDASWkAAPDaa9vWLBaL/quvvlp9/fXX6/l8vhZCbKSUu8taCLGy1i632+18tVrN27Y9tdYulVKrIAhWUsrVdrvdWGsbrXUjpdwSUXdycmLKsnSPHj3yH3/8sWeMEaEtFgB8RwhAAAAAAAAA/oTRWcsrRkTi5s2bYjqdSiGEDoIg9N5HjLGYiHLvfWatzbuuK9I0rfI8r2/fvj2q67qK47iw1mprbbC7OOd0GIY6TVM9GAzCMAylEAJtiQEA4LXX971r29bM5/NutVq1bdu2QoheCNEJITrOecc537Ztuzw9PT19/Pjx8WKxOOq67vTyjBAiWjjnVlLKVdd1GyLadl3X3bp1y37++efuShCCEAQAvhUCEAAAAAAAgEvBR1mWfH9/XxCRLIpCbjYbHcdxJISInXOJ9z7jnBfW2gERDTjngzzPR1VVjd59993JeDyukyQpvPfSe8+dc8J7z733QgghgiAQSikphOCcc/xNBgAArz3nnLfWuq7rbNd1zjlnOeeWMeY455Zzbr33ZrPZrI+Ojk6/+OKLw5OTk8PtdnvCGDtxzp0yxo455ydEtFAgITSHAAAgAElEQVRKLZxzK2PMhoi2o9Got9aaw8NDlySJG41G7pNPPnEIQgDg2+DDNgAAAAAAvO34hx9+yP/xH/+RPX78WCRJIowxQRRFARFpY0xMRAnnPLXW5s65nIhKKWUZBEGZpmlV1/WoLMvhzZs3R3Vdl0mSpIyxb8z18N4zxhidt+8gwt9kAADwZjgb1HE2r4O893Q1mHDOuaZpmpOTk8WTJ09OTk5OjhaLxXHTNCfOueO+748YYyec81Ol1JyIFudtszZxHG+jKGrbtu0Hg4E5ODiw7733nvm3f/s3T0RuNpt5QlssALgGyq0BAAAAAOBtxYiI/9M//ZPIskxKKYPbt28HURSFWuvEe58T0YAxVhPRyDk37rpuYq2d9H0/kVJOsiwb7+3tTabT6WQymdRFUeRRFEVSyoAxxtlznL82wg8AAHhTMCJ63tvepbc/YpxzppSSUkpJRKrrOrndboPtdqu895qI9O6aMaaFEIFzTnVdJ5RSvOs6obVmT58+ZXEc0y9+8Qv/7rvv0sOHD1/m/gPAKwoBCAAAAAAAvG0YEfF79+7xu3fvyiiK1K1bt1QQBKFSKpJSxkSUG2MG1tqKiEZENOGcT6SUEyHEhIjGSZKMiqIY7+/vj6fTaV2WZRFFUSilVJxzTgg4AAAAnsEYIyGE0Forzrm01qrNZiP7vg+stYEQItxdOOfae6+99wERSc45d84Jay13zvG+74lzTm3b0sHBARuNRvTo0SO89wLAM+TL3gAAAAAAAICfgveeffTRR/zu3bvs6OhIaK2lEEJGUaSklNpaG65Wq6ht22jX6soYU2qtyziO6yiKKillcb48jaIoLcsyK4oiz7IsSZIk3FV9vOx9BQAAeNUwxohzLpRSXEop+77neZ6LoigEEekwDEOlVMYYy5xzRdM0Wdd1p9bamDEWEpEmoqWUcs0Y2wghNm3bbq217a1bt7o8z810OnV1XdtPP/3UP3jwwBHaYgG89VABAgAAAAAAbzTvPbt79644ODjgYRhKznmQJElorY201knXdZn3vrDWDowxVd/3Q2PMuO/7sTFmHIbhtK7rvRs3buxPJpPpZDIZ1XU9GA6HxXA4TKuqipMk0UEQqCstrgAAAOBPLnphcc75+UwsoZQSaZoGZVmGdV3HWZbFWuu4bVvVtm2w2WwCY0zQ933gnNPW2sBaq40xylorxTmttRgOh+yv/uqvWJ7n7F/+5V/ovDUWQhCAtxgqQAAAAAAA4E3GHjx4wE9OTvh6vRZCCNn3ve66LoqiKOq6LpZSxtbalHOeMMYyIso55wURFd77QmtdZVk2HI1Go8FgkIdhGDvnJGNMCCFEGIZSKfWNgecAAADwfFJKkWUZBUHAjTGaiGLOuW2appnP5+vFYhEsl8vIORdxzmPGWOK9T40xS+/9UgixYIytmqZZZVm2Yow1jLFmsVjw6XTaN01DH3zwAXnv/dWB7ADw9kAAAgAAAAAAbyp2//59TkSiLEuxXC5lmqbBdruNhRBp3/fZ7pqIiiAI8izLijzPCyFEQURZ3/dZWZZ5VVVVnud1nudJFEWh9/5i2CvnnHHOUfEBAADwZxBCMM65kFJy770kooAx5oUQgfdeDQYDcs6pIAi0ECIhosxaWzRNs2jbdtF13amUci6ljPq+10EQLIMg4EopZq1lq9Vq91Lee+8QggC8nRCAAAAAAADAm4jdu3ePE5E4OTmRSZJIKaUiotB7nxBRYa0tnXMDIio452Ucx4O6rsvJZFLFcZwTUeKcC6MoSoqiSNM0TbTWoVIqeKl7BgAA8Aa41A7rmeVhGDJrLdV17cMwVGVZxkKIwjm36rpudXh4OD85OTndbreptTZRSkWc892gdLLWMmsty7LMCyH8o0eP/KeffkoIQQDeTghAAAAAAADgjTObzdgHH3zAPvvsM54kieScB0KIYL1eR1rrdL1el4yxkbV26JwrhRB1EAR1WZb1zZs3h3meZ0EQaOec5JyrIAiC82HpmKMIAADwIxJCiCiK9Gg0YmVZhsYYwzk3fd9vV6vVpm3bk8VicUpEqXMucc5FzrnAey+899Z774MgcIwxxzl38/ncvffee57OBqIjAAF4y6BMGwAAAAAA3hTs3r17/Fe/+hVfr9e7ig8thAiNMSFjLLbWpm3bVl3Xjfq+H0sph2EYVmmaDkejUXXr1q3q//2//1fmeR4HQaC89/zSvNbzma0Mf0cBAAD8SPw5d8afz/Bwbdv2q9Vq+9VXXy0eP368OD4+Pur7/sg5d0REh5zzA8bY0yAITrz3izAMl0KINWOsybKsLcuyj6LIPH361B0cHPh79+6hIgTgLYCzlwAAAAAA4E3AZrOZ+PnPfy6JaFfpERtjsrZtB9basuu6qm3bYdd1k67rJkQ0juN4VJbleDKZjKfTaTUcDgeDwSCL4zhSSmkppRRnEH4AAAD8BC61xuJCCHH+Viw558J7L733gnMuOOeCiHjXdbuLOK8CkdZaZa2V1lpBRFwpxZ1z7PDwkLVty8IwZF9++SW9++679Jvf/Ib+9V//9WXvNgD8SNACCwAAAAAAXmdsNpuxTz/9lFVVJZqmCaIoCvM8j51zSd/3uTGmsNYWRDTo+35gra36vi+FEKWUshwOh+U777xT13WdZlkWRlGk+NWG5AAAAPBScc55FEWyrutIa83DMORExNbrNW/bVnrvtfc+dM6lSqmTvu9TIooZY/Ou6xZt226iKNpwzlutdUdE7IMPPjBE5AitsQDeWDh7CQAAAAAAXjdsNpuxO3fusJOTE/748WOxWq1EXdeBEEKHYZhYazNr7S78qJVSZRiGlZSy9N5XbdtmnPO8LMv8nXfeyd95552iKIrofM4HZ4xxVHsAAAC8Os7bYnlrrWvbtp/P580XX3yxfPLkyWI+ny+IaCmlXAghTo0xJ8aYI2vtkRDiVGt9yjlfBkGw0lpvtNbb7XbbKaU6a62Josh++OGHjog82mIBvFlQAQIAAAAAAK+V+/fv85OTE75er4UxRmqtVZIkqm3bSCkVNU2TE1HR9/3AOVcqpUZa63o0Go3SNK2klKUxJvLeR1mWxaPRKM7zPE6SJMCQcwAAgFcTY4wJIdiuLaVzjtV1TUQk8jwPiSiTUg6MMYPtdpudnJzEfd9Hfd/HRBRyzuPzCpHVer3ehGHYWGsbpVT3/vvvd48ePbJ37tyx3nvMBgF4g+DDPQAAAAAAvDa89+zf//3fRVmW8osvvtBSyjAIgoiIEu99bowZGGOGXdcNd4POwzCcFEUxuXXr1v6NGzem0+l0PBwOi9FolA6Hw3gwGOgkSXaVH6j6AAAAeA1wzkkpxZMkUYPBQFdVFZdlmSRJor33arVa8aZpeN/3kjEmiUgyxoT3XjjnhHOOW2uZlJJtNhtaLpfsd7/7Hf33f/+3v3v3Lnv48OHL3kUA+AGgAgQAAAAAAF4HbDabsYcPH3IiUuv1OsiyLHTORdvtNiGiJAzDXClVKKWGnPPyfPD5IEmSejAY1FVVDeu6rtI0Tb334ny+KjsfsIrwAwAA4DXBGGNSShHHMdNaS+99wBhz1lrbNI3q+16sVivGGJPGmCgIglQplRFRaq09sdbOu64LiSho21Y550QQBE0URUREtLe35+7fv+8++ugjT2fzQVARAvCaQgUIAAAAAAC86thsNmN7e3sijmMhhNDz+Tyy1ibb7TbnnA+895XWepRl2WQ0Gt0simJ/MBjspWk6KstyWJZlNR6Pq6Io8jRNkzAMA621DIJASik555whAAEAAHg9sLOzGJiUkiulRBAEUp1jjO2qO0QQBCqO43AwGMRxHIdhGAbGGGWtlcYYIYQg7z0TQhBjzMdx7Pq+9+PxmL788kuKoogePXr0sncXAL4HVIAAAAAAAMCrjN27d4/v7e3xn/3sZ4KI5JdffhlKKZOu6wohRNn3fe29r4IgGOd5Prl58+atPM9rrXXR971mjGmlVJimaai1Vsg5AAAA3kyMMRYEgSyKIlFKCWNMSkStEKIzxixWq9Whc+6JMSYjosQ5p6WUmoiEtZY1TePiOPbGmP5nP/vZbrXuwYMHu9uoBAF4zeCTPwAAAAAAvGrYbDZjRMSJiN+5c0csl0sppQw458F8Ps+893nbtiXnvJZSjoMgGNV1PRmNRtPbt2/fzPO8CsMws9YKIhLnba521R6c8LcQAADAm8g755y11hljrHPOEpHlnNuu61bL5fL466+//vr09PTpYrF46r3/2nt/yBg7ZIwdE9EpY2zlnGsZY50Qonvy5Ilt29YeHx9bInKz2QwtsQBeI6gAAQAAAACAV8ZsNuPncz54nueiKAq5WCyUtVY750JrbdS27cBaO3DOVWEYjuI4nmZZNqnrelKW5ThJkmmSJLnWOnnZ+wMAAAA/KcY5F5xzoZRSl+8QQmhjjMyyjDvnpPdebTYbvt1uZdd1UgihiChgjIVCiA0RNcaYZjQa9UKIbjqdmvfee88QkT0PQQDgNYAZIAAAAAAA8Erw3rODgwOeJImKoiiIoihUSsXW2qxpmkHXdVXf96Ou6ybGmGnbttM0TfeGw+GNGzdu3JhMJtPhcFgnSZIqpQLOOU74AgAAgB1PRPx8/pcSQqimaXjTNGq1WgV930fW2tAYE3nvA865EkIIrbXw3oskSVjTNPSLX/zC7+/v08OHDxGCALwGEIAAAAAAAMDLxmazGf/f//1feXR0pKqq0t77iHMeE1FujCmdc7W1dtR13cQ5ty+E2IuiaFqW5d54PN7f29vbq+u6zvO8CIJACyEkY4y/7B0DAACAVwNjjM4rQwIhhGKMqaZphLU2cM6FURQlURRFWuv4vO2mdM4J77303nPvPWOMse126/I8p3v37tHdu3fZw4cPX/auAcAL4IwoAAAAAAB4aWazGafzWR9EJBljgTEm9N7H3vukaZqciAbe+8IYU1pra6VUrbWu0jQtB4NBVZblMM/zKkmSJAzD8OXuEQAAALyKGGNCSimklIH3XlhrRZZl/nwQeiql3AghBt77067rwu12G1hrhTEmYIxJKSX33jMhhBuNRuyzzz4zd+7ccffv37ePHj3yH3/8sWeMoSoE4BWDAAQAAAAAAF4GNpvN2AcffMA/+eQTGUWR6vs+EEJE3vuYiNK+7zPvfWGtray1Zd/3Vd/3VRzHw6qqqhs3bpRVVRXD4TCP4ziUUqLCHQAAAL6VlJJHUaTH43FRFEXQdV0mpey890tjzOnR0ZFyzsnVasWFEFpKqdq2lUII2XUd45zLd955pyUiQ0Tm17/+tX3w4IHz3juEIACvFgQgAAAAAADwU2JExO7du8c++OAD9tlnn8mqqgKlVGitjYgoMcZk1tpcCFFwzksp5dB7X0opKyllmWVZVVVVOZlMyqqqkjzPI6WU4pwjAAEAAIBvxTkXQRAEg8GAGWNC55zlnFtrbd62bdp1HTVNw7TWzDmnvfdB13WBlFLGcUzn4YhM07RtmqZbrVaGiMyDBw8IIQjAqwUBCAAAAAAA/FQYnc/7ICL+29/+ViRJEjjnwr7vUyFERkSFtbZwzg3CMKzSNK2jKBpxzsu+74u+7/OyLAej0SirqioviiKMokgxxl7yrgEAAMDrgnPOOOdSSinpbDg6EREZYyIppc7z3PZ9z733ar1ep23bJs652Fqrt9utiuN47r1fd1239t43jLG2KAo2n88JIQjAqwUBCAAAAAAA/GRmsxm/c+cOJyLRdZ1qmibknKeMsdJ7X3rva2NMxRirtNZ1XdejyWQyDoKgIKKk7/soDMMoy7IwjuNAKcUZ0g8AAAD48zCis8Hou9tERJxzFQRBlOd5LYQQSqnw+Pg4Ozo6ytq2Tb33sdZad10XSylPrbVKCCE457zrOiqKguq69g8ePCAicnQpXAGAlwMBCAAAAAAA/NjYbDZjdD7o/ODgQMZxLI0x2jmXWmsLxlhNRCPv/VgIUQdBUKdpOhoMBqPRaDRO0zTlnIfWWimEkEopobWWQgj+kvcNAAAA3hD8rCxEJ0lSSCkDxljUdV28Xq+Ttm1j731orVWMsdAYExCRcM5xxhjfbDYsz3N2dHRET548MbPZzBKRm81mnhCEALw0CEAAAAAAAODHwu7fv89HoxH7n//5H9G2rTTGBH3fB/P5XBtjYmttzhgbnAcfY6XUNEmSYZIkw6qq6qIo6izL6iRJ4vM2FYyI2A7nyD8AAADgh3H20YIzpZRgjCljjMqyTDZNE3jvVdd10hgj2rZV3nvFGJPeeyWlDIwxqmka5b3f/PVf/3X7+PFjc3p6an7zm9/Yg4MD/+jRI48wBOCnhyGBAAAAAADwY2Cz2UxYa2WSJMpaG/Z9HxNRdj7Lo+y6bmitHfd9P+m6bso534vjeG80Gk339/fH4/F4WFVVkWVZEgRBIKWU/E/YeesrtL8CAACAH8rFORZ0VhDCOedCKbWbFyKapuGbzUY2TaO6rgucc6rrusBaG/R9rzjnsu97Eccxz/Occc7Z8fExi+OYoiiiR48evex9BHirIAABAAAAAIAfEpvNZvyf//mf+Xm7KrXdbvVms4mstalzbmCtLTnnNWNszBibEtHEez9RSk3yPB/v7++P9vf36+FwWGRZFimlAiEEZn0AAADAT4YxRowxJqXcBSCi6zqxWCx40zTSGKMYYwFjLCCiwHsfcM4lEXGlFIuiiGmtqes6nmUZLRYL9nd/93d09+5d//DhQ1SBAPxEEIAAAAAAAMAPgdF5y6uDgwPZtq3abrfaWhtZa2PnXNb3/aDrukoIMdJaj8uy3Kuqaq8oir00TcdZlg2Hw2E9nU4H5+FHHATB5fADAQgAAAD8JM7Pu+BSSi6EEIwxbq1lXddxIYSMoijI8zyMoijQWgdEpJxz0lrLlVLMOSeMMdw5x/q+51prdnBwQO+8846/d+8e3b17lz18+PAl7yXAmw8BCAAAAAAAfF9sNpuxDz/8UMRxrIIgUEopTUSRtTZljGXGmEHXdZVzbqS1HhdFMZ1Opzen0+nN4XC4NxgM6qqqyuFwmNd1nRVFEWqtg/MDDgg/AAAA4Kd2aeQYZ0TEvPdcCMGTJAmKogjLsozjOA6DIAj6vpfWWmGM4UR00ULLGMPPV8KUUsQ592ma0vvvv0/vvvsuoRoE4MeFIegAAAAAAPC9zGYz9sEHH/DPPvtMOueU9z5o2zYUQsRCiNQYkzvnBoyxgTFmJIQYJ0kymUwmN8bj8SSO48F5GwkppVRhGCqttUTLKwAAAHgVMMZYEASiLEsdhqGw1sZEZDjntmma/OTkJN1sNmHbtoG1VlprlRAicM4F3ntFRPK8koSlaeqFENQ0DX3wwQfkvfeMMYQgAD8SVIAAAAAAAMBfzHvPiEj89re/VXmeB6enp7G1NpFSZt77gXOu7rpuJKUca62nVVXtjcfj/clksjedTvfKshxlWTaIoiiMoigMw1AppaQQ4uJsy5e9jwAAAPB2Y4wR55wJIbhSSmqtVRRFQRiGmjEmiUhYa4VSSqVpqqqqCvM8j6Io0kop4ZwTfd9zay03xpD33hMRKaX8f/3Xf3m0wwL48SAAAQAAAACAvwQjInb37l3OOZec82C5XIZCiNQ5lznnCmNMZa0dWWvHWutJmqbT8/BjMhwOx1VVlWma5lrrWJ4RYpd8oO0VAAAAvDouemEJIfj5ZxYphNhVrArGmIiiSKVpGhZFkWZZFoVhqPu+Z8YY3vc9CSEY59xJKT0ROaWU22w2/uDggD788ENCCALww0MAAgAAAAAAfy5GdNb6Skop+r5Xm80mlFLG1trcWjvw3tfOuZFzbmKMmUZRtFeW5f7t27f3p9PpeDweV1EUJUqpgHOOv0sAAADgdcWklFxrrZIkifI8T4uiKKMoSqWUcdu21HUdNU3jiYiEEC4IAieldFEU2TzPrdaaEIIA/DgwAwQAAAAAAL4rNpvNGJ0P9szzXLRtq5xzoTEm6bou55yX3vvSGFMzxkbnlR+jsiyHw+GwLstyWBRFFsdxfF7tgfADAAAAXlucc747ocN7HzLGLBG5vu+1MUZ67zd935u2bZ0QgnnvvbWWSSm5MYaHYciJqH/vvffM6empmc1mlojcbDbzRITZIADfEwIQAAAAAAD4NoyI2IcffsjpLPyQYRiq7XYbOOdCpVTsnMuJqCCi2ntfWWuHURSNsiybDAaDcVVV1XA4HAwGgyJJklBrrV/qHgEAAAD8ADjnnIi4EOKZ46zOOe69933fL7uu65um8Uop0fe9CIJAEVGgtQ6MMSoIgi0RbafTaae17suyNPfv37f37t1zGJAO8P0gAAEAAAAAgBeazWbszp077MmTJ+L4+FgRUcAYC6WUkXMu9d5nzrmi7/vSOVczxipjzDBJkmGWZeMbN26MhsNhURRFliSJllKi6gMAAADeaNZaYa0N2rZNN5tNtdlsnJSSK6WEMSYIgkB770NrrRZCLJVSa+fcpizLdrvdtmEY0oMHD4iI7MveF4DXGQIQAAAAAAB4HjabzdhXX30lbt++LZqmUWma6u12G1lrE+dcKoQYKKUGWZaVUsr6fPZH2XVdWZZlWVVVXdd1MRgMsjRNI6UUPz9TEgDeMM45cs5R3/dkrSXn3DP3n80Jfv7Xl3nvv9PjfmqXt4vom9t2+f6rj+WcE+eclFIkhCD8KgR4szHGOBEFQRCkSZKYqqpIKaWklAHnPDLGREQUGWMCa62WUioikkKIdZqmrCxL1jRN/5vf/IZ9+OGHFpUgAH+ZV+dTBAAAAAAAvEou5n3kea6klGq1WmnnXMw5T4go6/t+IKWs8zyvy7IcZlk2FkLU59UgWZqm2XA4LG7cuJHneR5FURS87J0CgB+PMYbatqXVakVd15Ex5pn7d2HBLhjYfX1dMPLnBA0/ZEDyotf13j+z7d77595/3bqklKS1piRJSGtNSqkfbLsB4NWz3W77xWLRfvnll6v5fL7ebrcrIcSacz733p82TXPYNM3Rdrs9EEIccc6PvfdzIcTSe79K07RxzrXHx8f9H//4R0OYCwLwF0EAAgAAAAAAV11Ufvz85z+XXdcF1towCIK467rMe5977wfOuVpKOZ5Op5ObN29O9/b2biRJUhJR6pwLhBA6jmOdpqnWWkspJSrQAd5gTdPQYrGgJ0+e0Hw+p6Zpngk5LocF1319+frq8l3Y8F3Ckd2yq4/7LnbPuRrS7JbttuPq45xzzwQg3vuLCpjdsjiOqSxLmkwmlOc5xXH8Z28fALw+jDG26zqzXC77rus6Y0wnhOitteuu6xZPnz49ODw8fHpycvI1Y+wpY+zwPAiZc85PGWNrrfVms9lsb9y40RGR+eSTT9zHH3/sUQ0C8N0hAAEAAAAAgAuz2Yx/+umn7O7du4KIZFEUwWaziZRSsbU2N8YUQoiBlLISQoySJJlOJpPJjRs39vb39/eSJBlIKUPnnBBCcM65UEoJfu5l7x8AnB2Qt9aSMeaibRXRNw/2f1vLqquP2Ww2dHp6Sl988QWdnp7SarW6CC2uBhzXLSM6axN13Wtffs7V6o/rqkG+SwBytZrj6vLrHr9b/+Vw42rocTn8uLy+JEloOBzS/v4+DQYDiuP4mde+WiHzou2++jwhBEkpSQjxSrUMA3ibee+dtdb3fe+cc9Za6zjnzhizbZpm/fXXXx8eHR0dHB0dfd113dO+758yxg699ydKqWOl1IKIVs65lZRyS0QdEdlHjx45OqsGcS/eAgAgwgwQAAAAAAA4w84v/O7du5yeDT/Svu8zzvmAiCrvfSWlHBZFMRkMBntVVU3yPB+naTqM4zhTSqHVFcArzFpLfd/TZrOhtm0vWlVdV5HxXb8mOgtA5vM5LZdLWi6XtF6vnxt4XFcN4r2/CECIng1DrqvIIHp+UPNdqz+eFz5cXu+LHrO7vnq5Wv1BdBaaaK1pPp8TY4y6rrt2P64LWq7b593rKKUoiiIKw5CCICAU2wG8GhhjXEpJUkpBRBc97/q+DzjnQVEUZIzhfd/zzWbD1+s177pOOOcUY0xwzqVzTsRx7Nu2pdFoRI8fPza//OUvzX/+53+S9x6VIADfAd4VAQAAAACA6KztFT86OhJ/8zd/I4hIbTabiHOeeO8L51zV9/3QOVcrpUZhGI6Gw+Hkxo0be2VZVlmWFVrrUAiBKg+AV5wxhjabDR0dHV20qiK6virjcgXH5QPz14UlXdfRdrulruuIMUZBEDzzmOdVdlz3es+7/zo/1DyQF80mubz9V/flRYHI5TCGc07b7ZaOj4+paZqL78/VsOby83df79Zzdbm1lpIkocFgQKPRiDjnCEAAXnGccxEEQVAURSaE4FJKcXh4KNq2lev1WltrYyIKiShkjCnvvc/znLquY1VVtVEUsV/+8pf04MED7713CEEAXgzvigAAAAAAb7eLeR/z+VzevHlTHh0dBWEYhn3fp0SUO+dqxthISjmRUo6SJBmVZTmu63o8Go3GRVFkYRiGUkrFGEMAAvAjsdZeXP500NwTMXYxEteTJ/acbte7A/ZN09BqtaSjoyM6Ojp6plUV5/yFlRpEZwfyry4jOjsgb4yhvu+JMfbMgfhvq8i4WuVxOUB4nucFH1eHkX8XV1tgvWg+ydVWXN+1dRURUd/3tFgsaL1ekxDi2tZbl+eKXF3vrsXW7rZzjrIsI2MMBUHwjeqT7xoIXQ53hBAXFwD44XHOmVJKJkmSSCklY0wYY3jTNLLv+7Bt29h7H/Z9r5VSous6HwQBC8NQGGMkEW3zPGdRFLGHDx8a771FCALwfAhAAAAAAADeXmw2mzEikvv7+zIMQ8U51+d/dCdEVBDRoOu6Eed8rLWepGk6KYpiXNf1sCzLOs/zMo7jWCmFvy0AfkTOOer7ntq2pa5rqe/7Px0Yv3ywnq6vtDj78mzZdtvQcrmk+XxO8/n8olXVdRUgu7Djahhl/rAAACAASURBVBhyeflVlyseLi+7bnj4bh3PCx2uc107rOe1q/pzXDcT5Nvagl3Xtup5GGNkjCFjzDcCm6vX11V77K4vD1zf3VZKUZIk5L2nruteOMfkRfstpaQwDCkMw4tADAB+WIwxLoTgQgjJOZfWWr7ZbGiz2QhrrVqv18F2uxXGGG6M8Uopa4yh9XotGWOqbVuptWZ5nlPf90REfjab+dls5ukiDgeAHfyRAgAAAADwdmL379/nRCT++Mc/qiRJguVyGRljYudcyhgr+r6vvPdl3/dDpdQojuPJdDqdTiaTUVVV5WAwSLXWgRACE3cBfmTOOeq6lo6Pj+j09JQ2mw05584O1tPu4Dsjzhh5fznw8N8INnZBymazIWvtxeDs6w7wX60Iua5d0/Puf95w8W87CH/dY14UoDxvXX+uq62mrgtm/pzZIi9qF3bdup7XZuxF7bA452StpfV6TQcHB7RcLklK+a1tta5ug3OOhBAURRFVVUV1XZMQAgEIwI+Mc8601qosy4RzzuI45oeHh/LJkyesbVtmrSV29stAhWEYKqVCxtiybVux3W6593772Wef0a9//Wt7584d99FHHzlCCALwDAQgAAAAAABvodlsxh49eiSSJFFCCG2tDcMwTDabTe6cK5xzNRENOee1UqpOkqTOsmwyGo1G0+m0HgwG2fkf4pKIcIQM4Hu4fDb/5RZHRM/O11iv13RyckIHBwe0Wq3ImH73oGeCirOuWLsD7bvKjj9VLDjnyFp7USmwO8h9eQD51QP1l+/bLXvR4HCi6wd479Z9XTBy3e3nzQ553hyO7+N51RxXQ5fLr335evd9vG5/nredL1p+df3XVajslm+324sQ47p1Xn7+5Z+xy9dCCErTlIiIoigiIQQppa4NvjjnF5fvM3cF4G23a4eVZVkopRRSSmGt5cvlkqy13HvP4ziWSqlAShl677X3Xp3/vvFSSvZ///d/lCRJ995775nzShAihCAAFxCAAAAAAAC8XRgR0d7enlgsFkoIoaWUcdd1sTEmd86VjLHKGDMRQkyCIBgmSVIWRVFNp9NhXddVWZZFmqaxlFLgwBfA92etJWMMNU1Dfd/T+Rm/RPSnA+S72RGnp3M6OTml1Wp58biz4g/2zdDj/KtdePHs7IpvVmtcd727vas2Ibo+8NhdXw49nHMXocDV2y+qJrlcgXH5vutu/1iufm+uqz55UbXLdw1orla2XBduXF7nda+3a3t13grn2u27rgLk8rJdeNL3PQVBQHEckzHm2jkuQggKgoDCMCSlFIauA3wPjDFSSnEpZXA+D4R3XcfW6zXXWivvfRhFUaaUSpxzSdM02jknu64jpRRprVmWZf78/yH79a9/TXfu3HGPHj3ys9ns+hQa4C2DdykAAAAAgLfHbuYHf/z4sSIiHUVRfD7vIzPGlMaYyhgzcs5NtNZ7cRyP9vb2BuPxeDAajYqqqpIwDAMhBGdIPwB+EMYY2mw2dHh4SKvVitq2vWg/dTk02G63tF6vrrStomdmgOzCj4sD6peWn61nN5+D6Oox+e9SuXD1gPzVKo+rB+YvD+S+HKJc97zd476tbdaPHYC8KNjY3f+8KosXhUQvun01CHnRuq+bUXLd9jwvMLn6uF04tQvK1us1PX36lObz+cWg9stzR7TWlGUZ1XVNSZIgAAH4fs4aFjJGQggWhqEcDAYRY4y6rlOc8zgIgoFzLm6aJjo6OtpVh9i2ba0/R0QkhGCr1Yru3r1rRqORm81mhLkgAETiZW8AAAAAAAD8+Lz37O7du/zg4EDmeS7DMNSc84iIUudc3vf9wFpbG2NGjLEx53wvTdPpYDAY37p1q97f3y/H43GWJEmolJKccwQgAJdcbmFlrb24fbmt1dX7vPdkraW2bWmxWNDXX39Nh4eHdHR0RKvV6pnLcrmkzWZDbduSc5aIzio7hBQkLrUj4lxctCW6CEkutcHaBSREf6pseNFciqsHynfLnhdCPK/t1eX1PS8oeN42XHXddv+Qvm39L9q+b7vvurDju6zveQHRLii7/JjLs1v4Mz8b37zsfk4uf72rKFmv17RcLmmxWNBisaD5fE6np6cXAZ3WmoIgICHEN37er7vsfvYvfw/wNgLwLMYYU0pxrbXKskzneR5mWZZorRURia7rrLXWGWOMlNIRkXfOeWOMN8b4JEm81pqOj4/p/fffp3fffZcePnz4sncL4KXCOw0AAAAAwJuNzWYz9tVXX4n9/X0xGo0kY0wtl8vIWpsTUdF1XWmtrYwxwyAIRkqpcRzHe2VZTkejUX379u10Op3GRVGEu8oPtjuSCgDkvSdjDLVtS13XfWOOx/Nma+xsNhs6PT2lL7/8kk5OTmiz2TxzcPry8/60Xn8p0Dg7vfdP91062393daUi4bqZEi+aR/GXVF08rxrhbfJDfg8u/7td39bsm69ztWrkun/jyy3Jdo/Zrf9yi6xdiJEkCQ2HQ9rf36fBYEBJkly7v8/7XkgpKQgCCoKApJQYtA7wJ/78/9zlwg7PGPPb7fZ0vV4fHB4efjmfz79aLBZf9H3/2Ht/YK09EkKcGGNWRVGsOeetUqrt+77/8MMPDRFZxhiqQOCthTpFAAAAAIA32C78+PnPfy4ZY5pzHrRtG3rvM+dcud1uh9ba2lo7dM4NgyAYnre9Gk8mk3o0GhXD4VAnSRKcz/x4O49iArzArorj9PSUFovFxUDqy2fmXz5gvXP5bPvNZkObzYaMMReVIVdbHf3pYPZZ+6qzZf7iNhEj7xzRbhkx8uSfCUGuC0J2nnfw+i9tOYVfFz/s9+BF7bGuLrv6us+rtLmuCmMX6F1+rLX2mfvW6zUdHh5S0zSktX7u61y+3gU3URRRURQ0GAwuAj4AIKKzAhC67rOW1jr23ld1XZPWOtBa65OTk3C9XsdN00RBEGgp5SljTHHON1JKEYbh9j/+4z9Y27ZEROan3x2AVwMCEAAAAACANxcjIp4kiey6LuCch0QUc85jIhpYa0dENLbWjs9vD6WUdZIk1Xg8rm7cuFHUdR1HUSSUUhh4Dm+ty2fCX3df3/e02Wzo5OSEnj59Suv1+iIAudpO6Wq7ol3YsasgITo7Q/5yQPHNdlHfHEx+ucX7WQjCyHl3EYIwYs+s87u0X4JX03XtsK5rY/a8CpHLj7/c1uzq8y+vcxdU7H6md4HfarW6mBNy+flX/89cDkDyPCdrLWmtL37Wn7efl7dl99oAbyPOeaC1zoQQSkqpvffBZrORTdNoIgqISHDOVdd1gnOuOOfs/Hm+aRrnvXfnVSD4pQ9vHQQgAAAAAABvoNlsxomI53muiqLQm80m4pynzrn0/7N3Lz1upNfdwP/nudSF91ux2ZJmxmPHhjGCERg2nFUwswiy8rb9Id4vMe2vM9oGyC6RtwGyCiIERhZjIL6M1TdeqlhVz+1dkEWxKUqaGeuu8wM4RbJJdnNEFruff51znHNd7/0ohJAZY06klNMoiiZJkmTj8XiYZVl/PB53h8Nh2uv1IiEENX9IM/ahacKJuq5hrd0dCb+/EGuMwXK5xHw+x2KxQJ7nB4PK6Vabn8O2RPvzQA4XrY8t+B4LY24tcjfnAzYVINhsjy0084Lyu+vYEPVDzwruvstj364+2mydc7datR0L1Q6DkBDCbl6IUgppmsJaC631rfsdPoaUEkopxHEMrTUPXWcfJCGEJKJYSqm996LT6aDf7wfvvZRSyu3nkyqKQiqlNBFRnucijmPSWtP//u//4t///d/d7373O//ll18GbonFPiT8qcEYY4wxxth75vz8XJyenkoA2jkXO+dSrXU7hNAvy7IvhBhYa8d1XZ845zKt9aTT6UxOTk5GWZb1syzrDofDtNVqaa019ydhH7T99lZFUaCu62cuBjftr4wxu2Bjv+Lj8H6NwwXs583cOJzbsX/d4flj92tw8PH+eFa7q+e5XT307Mc7PH8YujSB4OH3flYFiPceZVliuVzi8ePHtypIDueSNNdFUYRWq4XRaAQi4gCEfagEEQkiQhRFPk3T/mAwCEopkaapnM/noSgKUZal8N4r771I01QYYyhJEvr6668xHA7NZ599Zh88eOD2KkIYe+/xpwZjjDHGGGPvH4Ft+FGWZSuE0A4h9Ky1wxDCyBgzrqpq4pybWmsnSqlxv98ffvLJJ4PZbNYdjUatVquloiji8IN98Jp5B3/9619xfX2NPM+fam3VzEWoqgrWbtqsCyGeCj8OQw4At65rrj82n6O57f72WGDyrLkeHHh8OJ712jp2mxe10zp2GcCtmTbPC+WabdNqi4h2FVN1XT9VQdIEH83Q9RAC2u02+v0+tNbQWiNJku//P4ex94CUUqVp2hZCqDiOdRzHuqoqX5YlWWtFCEGFEISUUjQVvFrrIKWkH/7wh0jTFA8ePAAA9/zvxNj7gQMQxhhjjDHG3g90fn5O2La9yvM8UUq1iKhrjOl77wdxHGdpmk7SND3x3o+ttZOyLAedTqc/Ho/7s9msMx6P036/H0kpue0Ve+8552CMQV3Xu/ZTwO0F36ayoxlwvlwunxpuDuDW4u1hONJ8/XlzGhrHZjIcOmw5dHj94XXsw/Ssf/vnVQwdCz9eNGfk8Hb7l/dn3+wHJlVVwRize4z9io/DEKSua3jv0ev1AABVVe3eX0qpXTDClSHsQyGEEEqpSAihms+gwWBgiEgIIbS1NrbWqqqqlNZaSCmFc47W67UEIJbLZd3pdMz290Z/fn7u3+gTYuwV4yO6GGOMMcYYe7cRAHF2diastbLb7aptj+h2CKHnve8bY0YhhHG3250Nh8M70+n07mg0mg2Hw5N+vz/Msqw3mUza0+m01ev1ojRNlRCCiFdO2XsshIC6rpHn+S7caOZ3FEWx2zbX39zcIM/z3WLs/twO59ytBdz9VkGH3/PY4nMTehxe/6zLAG6FLM/6fowdc+y187zX7LEQ40WeN29mP+ho5uo869S8N4QQkFLCGIOqqrBcLlEUxS4MaYIQxj4QtA07JG2I7RVSCCEBiKYqEQCklEEp5Z1zYfveCmVZ4uOPPw5//OMf8cUXX+Dhw4fcDou9tzgeZ4wxxhhj7B12fn5On332GT169Ej2ej2plNLe+8Q513bO9ZxzQ+/92HufxXF8OhqN7n700Uf3Wq3WWErZc85pKaXWWutut6ujKBIv/q6MvfuaI8sXiwX+/Oc/78KNpqqjOarWe7+rEiGio4usL6rEeN7XQwgQQtwKQb7P0GrGXoX91+qx1+ixipFmvsjhe+CwKgTAbv7H/u32A5Lmseq6xuXlJZbL5W6QehzHaLfbuzkhSZJwEMg+OFJKmWz6wo211lEURbH3XuV5TtZaEkI0n18+iiIYYxBFUWi327i6ugq/+tWv8B//8R8AELYnxt47XAHCGGOMMcbYu4maYeeXl5daCBEZY5I4jlsAuuv1euS9H2utp61W66Tb7Z6enJzcnU6np1mWzXq93qjb7fbSNE1arVbUzPwQ29KPN/3kGPtbNJUZdV2jqqpbp7quUdf1bhDz9fU1Li4uMJ/Pd0POy7K8dR9jzFMtso4NNT/WIujw5zo24+PY5cPHY+xNORx+/rzbvehxDrfH3ktN+NjMB2kqT5rQsixLrNfr3fsyiiJIKUFEu/f4/vt3vV6jLEuUZblrd3f4vBh7lxGRkFIqIpJEJK21FDZvVlJK0TaYDNZa2lYrklKKpNwsCyulws9//nOuAmHvLa4AYYwxxhhj7B10fn5Of/rTnyQA3e/3IyJK0jRNjDFt51zPez/x3mftdvtkMBjMRqPRaZZlp+PxOOt0OqNWq9XWWvMkWfZeasKP1Wq1CzOA2wuv3nsURbFrbVUUBay1z2wNdDjD4Nh2fwYI8OwQ5NjXDucnMPY2et5r89vMrTkWFh4byN5UeTQVIk3LusP2Wd57XF1dAQDW6/VTj3NYvRJFEVqtFrrdLpIk2YUtjL2rtu2vhBBCYdMWlay1AQCklFFRFKooClVVlQQQSSmjEEJzkkQk2+02ffLJJ/jqq6/Cb37zGw+uBGHvGQ5AGGOMMcYYe/cQANFut1W/348ApEqptve+S0Q9Y8zQWjsloiyKotloNLrz8ccf3x0Oh1m32+0lSZJu/1Bm7L3knENZlri+vsb19TWKogBwe6E1hABjDMqyhDFmN0fgeY95rErjWW1+GGO3HRuUDjz7PXRsAPvh14wxmM/nqOsaWuujc0b2t51OB6PRCEopnhvC3jtCCBnHcdzr9fpSShHHcfz48WNRFIVar9dSShkppSIAkfdee++FUkoAwGg08nfv3nXn5+fh/PycP8TYe4X/6GGMMcYYY+zdQfuVH9PpNM7zvKW17njvewD6UsqhlHLc7/dPtNYnk8nkZDQazQaDwbTf7/fjOG5JKZXgw17ZO2p/cHIzIwC4vZjaDDefz+e4ubnBarU6Ouh5f9jy4RyO5rGa79l40WyDw7ZWjLEnntf6rfGiaqjDVnNNiLn/sXYYfjSnZpZPq9VCCAHW2qfez80MoCYkadoEMfa2E0IQAJ0kidh+3smyLF1ZlmStJWutAqCstco5J4mIQghie7/wxz/+Eb/61a/q8/NzB8BvgxAOQ9g7j/fijDHGGGOMvQNCCHT//n3x+PFjNZvNIiJK67puEVHPWtsPIYycc5MQwjSO45N+v39nPB7PptPpyWQyycbj8ajdbne01jHP+WDvMmvtLuBoWlc1MwHW6zWqqsJqtdrN91gsFiiKAsaYW6e6rndByr5nvTWahdoXVXfw/A7Gnu/YMHTg9nvncN5Oc76ZC9JcBjZBprUW1trdDJDmPX54AjazRaSUu1Z56/UaRVEgz/Nd27wmUJFScgDC3hm07YUlpZRCCAlAOudECEF67yUAYa0V1loyxpCU0jvnIKUMROSb94lSij7++GMAwKNHj97oc2LsZeAKEMYYY4wxxt5yIQR68OCBwOYApoiIEiLqCCG6IYSB937ovR+HEMZCiCxN0+npxnQ4HA673W43SZKEiHgVh73zjDFYLpd4/Pgx8jxHWZZPDVX23sMYc2uux/7Xm/P7gcbhUeeH1SDHqkCODT3n4IOxFzt8Dx2+n57XLutYNVdjvwpk/3vsD1JfLpcIIeDq6gpKqaeqROI4RrfbxWw2gxACURS9qv8NjL0yQgiRJIkejUbdJElkq9VS33zzjarrWhdFoZ1zkfdeRlGkrbVKKSXTNNVSStXr9YrFYlGfnZ3VZ2dn+M1vfhMA+Bd+U8beUvwHEGOMMcYYY2+x8/Nz8fjxY/Ho0SNZFIUmokRK2RFC9L33Q+fc2Hs/UUpN0zQ96Xa708lkcnJ6ejo7OTmZ9Pv9fqvVammtNVd+sHdJ0+rKWnurcqNpbXVxcYH5fI7FYrGr/liv1yjLEkVR7I4EPxxMfqzlzrG2VvuOhRs864Oxv82L2lt9l6/vhyLHrgewC0EA7KpFmsqPZrtcLneVYVEUIY7jWxUg3D2SvSu2r32hlJJCCElEctsGi6y1Apt5ctubEjWXt6Gg996HoijCxcUF/uEf/gEPHz7kDzz2zuIAhDHGGGOMsbcX/b//9//E9fW1EEIoY0ycJEkaQugaY4bGmLFzbqK1zqIomvX7/ZPRaHSSZVl2cnIyGY1Gg06n046iKOLwg71Lmt78dV2jKIpdsNG0t1osFri+vsZqtdpVeTQtrZqgxFp7dEbI4fd5VhXIscuMsVfjWRUdz7rt/vbw/LPaZ+1XiDX7irquUZblbv9SVdWuLV4URbsZIE0VCbfDYu+K/XZYcvPCFc45sQ0/BBHR9nOSvPckhCApZRBCBCmlIyKvtXbj8TgMh8Nw//798PDhwzf9tBj7XnjPzRhjjDHG2NuJzs7OxJ07d0Se50oppb33qfe+Y4wZGWMmADLvfSalPBkOh7O7d++e3Lt3b3p6ejoaDofdVqsVK6UkEfEhq+yd0gwyXy6XuLi4wNXVNW5u5lgul1gsllitVqiqEs65W0OLDxdRD8ONJgxpqkIOqz6OBSKcGzL29jhWvfVtbn9YIbK/z2jON/M+lFK7ahHnHLz3EEJAaw2tNe8T2Dtp+1oXcRxLrbUkIlFVFdV1Lbz3QmtNzSwQIYQNIXgALk3TMJlMQlEU+OUvfxm4EoS9izgAYYwxxhhj7O1DZ2dn4v79+/Ivf/lLtF6vYwCtEEIvhDAwxkyI6ERKOY3jeNbr9Wbj8fh0G36Mh8Nhr91up0opbnvF3jpNEPGsqo3mcp7nuLm5weXlJW5urrFYLHetaqqqhDH2Vn//YwOVm8XPJvBort+/zbN+RoDneTD2tnnee/LYXJHDr+/vL/bDj8NTU4XWtMNSSu2CkcO2fE2rPefcc+eTMPYmCSFIay2jKFJKKRlCEHVdUwhBElEzND0454K11gkhgtbaA0Ce5+h2uwFA+OUvf8ntsNg7h4egM8YYY4wx9pY5OzsT//iP/6iurq70aDSKvfcJEbWJqO+9H4UQxlLKSRRF006nM+33+9MsyybD4XDY7/d7nU4nldyng72lmvBjXZabAMRYAADR7UHHeZ5jsVhgPp8jz3PUtdlbuLzdBudY66pjFR7HHLueFy8Ze/c8K+Q8FkjsX7cfmjRVYiEElGW5C0+TJIGUctceq9nvNPdVSiGOYyRJAq01t8pibxUioqYVVlMZvG0xGQCIoiiEMUZYay0R2RBCZa311lofRVHTMgvD4TD85Cc/4YHo7J3DAQhjjDHGGGNvDzo/PycAUkqpO51OUpZl23vfATAEMLTWjo0x0yiKTtrt9vTu3bsnWZZlk8lkOBgMWlEUaa74YG8z5xzWZYmrq+vNAPOi2IUazYDhpgVWM8zcOb8XdASEgKcWL/fbWh22seJZHox9mI6FHM3l/euPBaZCCHjvUVUVrq+vUdc1Li8vb92mCUzSNMVgMECWZbtWWoy9jYQQFEWR7Pf7SQihn6apuLm5oYuLC1qv13YbengAUikl67qOpJQ6TVOhtQ4AwrY9Vti+p/gDlr31eI/MGGOMMcbY24HOzs7E3//938sQQmStTbfhRw/AkIiyEMJUCHEihDjpdruz0Wg0vXfvXnZ6ejoaj8f9VqsVR1Ekue0VextsFgc3PfSds7uh5GVZIs8LPL54jMvLS1xeXWGV58jzHHlebLebVlfltkrkyeLk0zM9joUd3vujlSGMMXboRdVhTTuszb4rx2q1wnK5xHK5xHy+mU1kzKZCLY5jSCl380Occ7uWWfut+LhNFnuTiIiUUiKKIqmUEt57WZYlbdu5EbAJSrbnSUoJa20QQrjFYuGJyP/3f/83FUVBjx49esPPhrEX4woQxhhjjDHG3gJfffWV+Mtf/qLSNFUA0qIoOkqprrV26JwbV1V1GkVRFsdxliRJNplMplmWjbeVH71ut9vi3IO9Tbz3MMZivV7DWrM7UrqqKqxWOW5u5ri5vsFqtQIASNkMJd7cfxNgHFZw3A469tvWHPb958oPxtgx+1UfzeXGYWsrALsg49hcoaYlljEGUkokSQJrLaIouvXYIQRIKRFFEVqtFqIoglK8JMdePyKClFIIIYSUUgEQxhhRFIUAEPI8J2MMOeek915qrRU2lcnknHO9Xi8sl8uwWq3s2dmZPTs7w6NHj8L5+Tm3xWJvLa4AYYwxxhhj7A0KIdD5+bn4t3/7N91ut6PlcpkWRdEty3IAYGiMmTjnMufcLEmSk16vd3Lnzp2Tu3fvTk5PTwej0ajdarVirbXaph/NibE3qq4NiqLYVHlcXuHq6hKLxZMjplerFcqygnPuqeADwK7i48l5PHX52KyPxuEiJmOMHc4E+TYh6f68ocPrmsdo2vc555DnOebzOa6urnB1dbXdB15iuVyirmsopaC1htb6ZT41xr4twqYIhLA5AyEElFJSa01KKaqqiowxZIwBAHLOkZQyeO+9tRZVVSFNU/LeU5qm4e/+7u/w6aef8nB09tbiuJkxxhhjjLE3JIRAAOjhw4diMBiom5ubxDnXds71rLVDIcTQe58ByLTWJ2maTnu9XnZycjK5c+fOcDgctuM41tvw400/HcYAPDky2pgaeZ7j8vIS8/kc62INEk+Orq7rTVXI7cHmTx6n6b8PbK7fH07cOFYFcng0N2OMNZ4XfBxWhuzfXgixCzqafVizj2pORVHAWnsrDGkqR7z3aLVaGAwGSJIEURRBa723/+N9FXv9hBDQWotOpxNFUSTjOPZCCBRFEZr2k9ZaIYSgsiwRx7FtXqtFUUghBKVpGtbrdfOQT45cYOwtwhUgjDHGGGOMvQH74cd//dd/SWttslqt2gD6dV2PvPcT59xEKZUlSXLS7XZnk8kky7Jscnp6OhiPx91Op9NSSqntzA+AKz/YG9b0uy/LEqvVCovFApcXl1jMF8jzHFVdwZpNP3y3DUqeHF3dPMrtocSHbWc2tz3evoYxxr6P/dkczfaw8uNZlSD7IawxBmVZ3jqt12uUZQnnHIhoNyekGZTeHIHP2JtARCSlbNphUQiBnHMEQDjnKIQgQgi0Df28UgpRFAUhRBBCOO+9F0KEXq8X7t+/H7gKhL2NuAKEMcYYY4yx149++9vf0unpqYyiSA4GA3l5eZl47zve+yGAiff+xHufKaWm/X5/eufOndlkMhkNN1pJksRKKT6gib1VnHMo1yUWyyUWiwXm8zmqqoL3DkAAAiEgbKK6vSWSwzkf+wFI8/V9XOXBGHuZDkON/XD2sDLksIXWYTus/fs3FR5NZdx6vcbFxQWcc6jrGsPhEL1ej+eBsDdl1wlLKYU0TbX3PgWAOI5lHMfi8vJSF0WhjDFKa40QgnTOCSISIQSvlPJaa3/v3j0PwIUQiIg4BGFvFd7DMsYYY4wx9nrR+fk5ff755+Lrr7+WRVEoItJlWaYAugCGIYSJEGJKRNNWq5UNBoPpnTt3JlmW9fv9Sk1IYwAAIABJREFUfmfb9ooPF2Vv1H5Lqmaxr643ba+ur66wWCyxXC5hnQUJgSiKNrfduw+2rWGOz/vAU5d5pgdj7HU43M/s7+cO54gcu31zn2bbtOhzzuH6+hrGGBhjIIRAHMe7eSCHFSi8v2Ovk1JKttvteDsPRBKRKMtS1nUtqqoSzjlf1zU11R9EVAshauec8967s7Mz++DBA4QQPIcg7G3CAQhjjDHGGGOv0fn5OQFQv//971VRFJExJtFaJ9gEHyPn3ERKmSVJMk2SZDoejyfT6XQ0Ho97/X6/3el0EiEECSF4VYS9MdbaJ62snIMPm8W9cl1isVjswo91ud4tAu7P9MCutZVH0zL8WcPM9/FiIGPsTThW6XF43X4bq8NZImEv7F2v17v7tlotaK2xHTYNANi2GEIURVBK8X6PvTZCCKG1Jiml9N6TMQZFUSCEACkliMgC8MYYR0Q2iqK6rmsHgNI0DY8ePQo///nPzYMHDyyA5gOesTeOS+YZY4wxxhh7fegnP/mJms1mkRAitdZ2jDG9EMLAOTc1xpzUdT2L43g2GAxm0+l0OpvNxlmWDcbjcafdbsdxHOvNyA9eEWFvhvcept4siszncywWC6xWK+R5juW29dVyuURZlTCmhvebSg/gyaLhphKEZ3gwxt4Nxz5yD1tlHdseng8hwDkH4EmoUtc11us1bm5usFqtUJYlhBCQUkIpxfNB2GtDW2LzoqPtSUophVKKnHPBWouqqhA2PBEFIoK1FiEEv1qtwscff+yn02l4+PDhG35GjG1wAMIYY4wxxtjrQWdnZ+LnP/+5Xq1Wife+Q0R97/0whJA552bGmJm19rTdbs+yLJv94Ac/yE5PT4eTyaTX6XSiZuD5m34i7MMWQkBZlpjP5/jmm29weXmJm5ubTfCxWCLPc5TVGtYaeL+p8vD+yWk/BPHhSRutpkUMY4y9K/ZDkMOZRYdtsw7DXu896rrGarXCfD7H1dUV5vM56rqGUgpJkiCOYw5A2BujlBJJksg4jqXWWhRFQev1er+KKUgpm7DOK6V8CMFfXV35H/3oR/7TTz8FD0VnbwNugcUYY4wxxtirRefn5/SnP/1J/vSnP1VVVSVKqXZd130AoxDCiIjGSqlZHMcnSqnTyWSSTafTcZZl/cFg0Ol0OolSioiIV0HYK+W9h3MOVVXDWgNrLQDCpuMagWhzmzzPcXNzg/l8jtVqBWvtNrwIcM7DB38r1NjM+8Cm6iPgqQoQnu3BGHtXPWsI+v51xwaoO+ewXq8BYBcQSylhrd3NBWnCEACQUkJrjTiOuTKEvXJSSiIiuT32JhBRyPPcEZFXSsE5FwC4/fZtIYSwrQQJAHB2dmY+//xz/7vf/c6fn58/GfbF2GvGAQhjjDHGGGOvDp2fn9Pp6akEoBeLRaSUallru865gZRyaK2dhBCyOI5P+v3+yWAwmGZZNjo5Oel3u912q9WKoiji39vZa+GcQ1lWWMwXm0qOstws2AkBIQhCCIQQUFWbWR9FUaCqK1hrIfYW/fzeIuCtEARA8HsLg3jx3A/GGHvb7Ye4x/ZphwPUm+ucc7cq5Ky1yPMc19fXAIBWq7ULOpIkQafTQb/fv3U9Y68CEZGUkqSUSNNUe+/DaDTyUkqvtUae53a9Xtd1XbttKywfQrBE5IQQTkoZsGmhZX/961+7zz77zP/mN7/huSDsjeA/pBhjjDHGGHtFtgPPxZ///Gcdx3HsvU+IqA2gR0SDuq5HIYSx9z6Lomg6Go2mH330UdZUfrRarUgpxW1r2WtjrUNZlnh88RiXF5dYLpcgQZBSQggJKcV2mLlDXdeoTf0k2Ng+xm7btLnaa2112CKGMcbeBy+qYDs2C6S5brNP3QQgAGCMwfX1NYqigJQS3nsIIdDpdDCdTm8NSGfsdZBSilarpcfjcTtNU6RpSo8fPzZVVdV1XTvvvQPgvPdGa223J//Xv/6V1ut1Hcex+eEPf2i3QcmbfjrsA8R7S8YYY4wxxl4NsT2pJEk0EaXW2i4R9a21I+fcRGudxXE8jaJoOp1OJ1mWjbIs6w0Gg3a73U6UUkJKyX8pslfK+wDvHax1yPN8N8ujGXBOQmzbrTRBiAAQdu2ymkW7WwPOv0UvfF4EYYy9jw73b8f2d0013X4I0tw2hLAJmOsaAG4FI3Eco9PpQEqJEAKUUnv7ZcZeDSGE0Fqj3W4LKaUXQvi6rmtjTB1C8FvBWmullC6E4Lfhnez3+0We5wSgmQfiwFUg7DXjo8kYY4wxxhh7+ejs7ExIKdV4PI6cc2kIoee9HzrnJnVdTwGcpml6Mh6PZycnJ6enp6fT6XQ6zLKs2+l0kiRJIiGEIF4lZq9YM/Mjz3PM53PMb+a4urrGcrlCWZUI3sM5C+88rLNwzsFaC+/dU2HGseDjGH5ZM8beV4f7t/3Lz/ra/rapnGv2tdZu9rvAJijZf4wm/JCSl/fYq0MbojkwZ/vrKRGRkJthIcI5R977QLRplymEgNYaUkqvlArz+TxYa/2Pf/xjz4PR2evGFSCMMcYYY4y9ZNuh52I8Hkuttfbep865XghhZIzJQghTACdJkpyMRqOTTz755CTLsmGv12unaRpLXslgr5G1DlVV4eb6BpeXV5jP56iqEkIQkjjeLLYRDkKOgBCeBBzNEcpPvs5trhhj7NDh/nE/zGiqOPbDkP3WWESEoijwzTffwBgDY8yuAkRr/TqfBvuASSlFkiTRYDDoKqUoSRJ9cXFB1lpaLpe+qW7y3lMIgcqydN77EEWRW6/XFk8qQPiXBPbacADCGGOMMcbYy0NnZ2fi8vJS/fjHP1ZSyrgoijYR9ay1AwBjrXWWJMk0SZKTLMumk8lkMp1OB4PBoJOmaayUktz2ir0KzYDd/aG7AFBVNVarFW62La9Wq9XuaGOlN38yEu23uNo83mF7qwYHH4wx9mz7VXPHquH2j4FoFpOb+xhjYK0F0aYlYZqm8N7DGLO7fXPkPVeGsFdBCEFSStVqtWhb7SGqqnJ1XQfnnN8OP99VLymlXFVV2IYg4Z//+Z/D559/ji+++MIREf/CwF4LDkAYY4wxxhh7Oejs7EzMZjOVpmlkjImqqmoJIbre+4FzbkRE4yRJsk6nMx0MBtMsy7LJZDLs9XrdTqeTaD6Ek71Czm0Gl+d5AWPqXchR1zWKvNiFH2W5BpHYDuvdf4SwvS7A+6fDDw4+GGPsxQ7ngxy7/tjtQgi7ELup+kiSZDcbpJkJEkUROp0OkiThAIS9CkJKiW21MoUQRK/X8845EFGoqio450Jd14GIgrXWeO+D1tprrV1VVT6OYzx8+BAhBA5B2GvBAQhjjDHGGGMvwdnZmbh//75M0zSy1raccy2tdW8bfkyttTOl1Kzdbp/cvXt39tFHH50Mh8Nhv99vt1qtSErJE0zZK2WMwXK5xF//+hh5nqOqKhBtK0OMRVGsYUy9XZDbtrRq2lxt+9I3w8+/7awPxhhj3473fhsy356pdDhDhIhQ1zUWiwWcc7tqD+89kiRBt9vF3bt3uTUWe+W27bD0aDTqJEkiWq2WvLq6EtfX16IoConN/PQQRZH03gtjDA0GA2q1WlRVVdMGy73hp8E+AByAMMYYY4wx9reh8/NzAiABRM65RAjRllJ2jTFDIhorpaa9Xm/aarWm4/F4mmXZeDqdDvr9fidJkkQpJYmIAxD2UuwPz92fzVEUmyqPm5sbLJdLrNdrSLlpr4LQtKtwT2Z8bO+3udjM/Qjc8ooxxl6BZwUfh1UiTdhR108q+YBNlV+r1YIxBp1OZ3e75n5N26xmbghjf6vtYHS0Wq14MwudYK11xhjvnPPGGA/AeO99XddBCOGrqvLe+2Ct9Q8fPsRXX32Fs7Mzz5Ug7FXiPR5jjDHGGGPfnzg7OxOPHz9Wn376qSaixHvfBtDz3g+89xMhRBbH8Wmv15uNRqNZlmXT2Ww2mkwmg3a73YrjWAshBB1rBM7Yd9S0SKmqCqvVCkVRoCgKlGWJ5XKJ+XyB6+srLJebrxljUNcG1jVhyZO5pE+CjifhR3P9/vdjjDH2cjSzPr7NrwTNjIW6rlGWJbZzFkBE0Frv5j4VRYGqqmCM2QUoSvHx0OxvR0QkhBByC4Dw3pNzToQQCEDw3jvnXAAQlFIegJdSOueci+PYL5dL/+jRI9y/f58ePnz4Zp8Qe2/xHo8xxhhjjLHvjgDQF198IWazmfz444+VMSbx3restV0AAwAja+1ESjntdrsnd+/ePZ1Op7PhcDju9XrdOI4jHnbOXrYQAqqqwmKxwMXFBdbrAtY6CCFgrcV6vUZd1wACpBTbWR9P7rtf3UG7tlfHgw4OPxhj7OVq9rv71R/7++LmNsBmWLr3HkKIW/erqgqPHz/GcrmE1hohBGit0Wq1kGUZRqMRoij6ViELY9+WEIKSJFG9Xq8tpUSr1Qrz+dxdXFzUeZ57a60nIu+cc9Zap7W2eZ6HLMsCAHt6eupCCA4AuBqEvWwcgDDGGGOMMfbd0RdffCF+9rOfyfF4rI0xcRN+CCH6IYSxUipLkuSk2+2ejkaj0+l0Ojs9PZ12u91ekiSx1lpx2yv2sjRtr4wxKIoC19fXuLh4jNVqBWMMhJC721lrEUK4tWj2rMd8XisWxhhjL9/hfvkw/NgPSJpWVk14TUQwxmCxWGC5XALYtMaK4xidTmfXAqupMtlvjdWcGPs+iIiUUqrT6ZDWWsRxDCLyZVla7z2MMQAA55xTSjnvvUmSJBBRiKKo+tnPfmb+8z//E//yL//iAPAvG+yl4gCEMcYYY4yx74bOzs4IgPj4449Vu93WZVkmZVm2hRBda+0gjuNhHMeTbrc7HQwGJ5PJ5GRb+dHvdDotKSX/Hs5emhACnHOo63o352O5XGCxWNwKQKSUu0WzJvw4fJz9ChBudcUYY2+fZt99GJQ0Mz+axWbn3C4cj6II1lq0221EUbRrldVUhyRJgjRNdy2yGPuuiIjkHiFEqOva9Xo9AyCUZRm2s0Fq51wNoIrj2LVaLQcgWGuxXC43U8dCCFwFwl4m/sOLMcYYY4yx7+j+/fs0n89lnudaKZWEENpRFHVDCAPv/VAplfV6velHH310mmXZ6WAwmG7bXmmu+mAvW7PYtVgscHV1hfl8jsVisW19JaE13Vowa+4D3A49OORgjLG32371x/6A88OvNSG3c24XalhrcXNzA2stLi8vdyFImqYYjUaYTCYQQnAAwv5mRERaa93tdttE5Nvttlgul7i6uvJVVVXOuTqKosp776y1TggRtnNp/K9//Wv329/+lsBVIOwl4gCEMcYYY4yx7+Crr74Sjx49Uv1+X2utYwBpCKHrnBuEEEbW2rGUchzHcTYcDqeTySQbDAbDOI4jpZTmYefsb9Ec3du0pyKi3ZDb+XyOy8tLLBYLVFW1W/jab5FyuH1e1QdjjLG3y/6vEE0Fx7H5IPvnm88A5xxWqxXKsgSAXQDS6XQQQkCaprvh6FJKDkLY97atBlFpmqZSShFFEQkhfFmWLoRQmU0/rCYAsUIIL4QIcRz7uq7d559/HrAJQPiXEvZScHM/xhhjjDHGvh06OzuTRKRHo1EkhEhCCJ0QQg/AuK7rzFqbWWuncRzPut3u9M6dO7Msyya9Xq+ntdZSSrFdkOAQhH1nzjk451CWJdbrNYqiQFmWKMsSy+US19fXuLq6QlEU20HnxxfD9sMO59zu681iGGOMsXdHE4bvt8RqKkCaU3M7Y8xTnyHOOQghEEXRLvRo7s8hCPs+tq8dIYRQ25l3EoDw3hMRhW2lkQ8hBGOMX6/XsNbuWl+122384he/QJqm9OjRozf9dNh7gAMQxhhjjDHGXozOz8/ldDrVSZLEzrmW1rptre0754ZVVZ0YY7LmpJSatNvt0XQ6HfT7/U673Y63ra8IHH6w78lai7IscXNzg8vLS1xdXWG5XGKxWGA+n2O5XGK9XsMYc3R+x+F2vwc8AA4/GGPsHXMYch/OBzmcE3LYDnH/Pt57WGsBAFprKKV4KDr7vgibQpDdC7QZkh5FERERbcM4qqrKe+/Ddl5NkFKG9XqNfr8ffvSjH4X79++Hhw8fciUI+5twCyzGGGOMMcZe4OzsTGDzu3OUJElS13XbGNP13g9CCBOl1JSIplLKjIhGSqkhEXVDCEkIQW4OaOPFZfb9NO2ujDEoigI3Nze4urrCarXaLXA1c0CMMU/N92jOP2u73zeeMcbYu2W/FdaxfflhKCKl3H1OAJvPmDzP4ZxDXdcIISCO4107rMO5IvuhCWPfAkkpVZIkLSml1loHIkJZlr6qKqzXayelDNZaaK1DnudBa03dbjeMx+OQZZkH4F/4XRh7Dg5AGGOMMcYYezYCgNlspgBE7XY7Wa/XbSll1zk3iON4rLWettvtUyI68d5P6rruJ0nSHwwG3SRJYsmHT7K/QXNEbl3XKIoCq9VqN+R8uVwC2CxKHZvlsX/k77PmfHD4wRhj775jLQ6b7bF9fBNmNJ8NxphdK6w4jtFutxFCgNZ6F5porZEkCbTWXBnCvrVtOyxJREJKqQFY55zrdDoeQAghuLquXQghrNfrkCRJ2IwIgV8ul/7evXsuhOC2j8WVIOx74QCEMcYYY4yx4+js7EwMh0MxHo91FEVxWZZtIUTPWjsCMGq327PhcHh6586dT+I4nimlRnVdp0qpNEmSdDgcxnEcS15gZt+Xcw5VVWG+bXO1mM+R5/nuKN2AgOC36wHbzX4FSFMdcmy4OYcfjDH2fjlsa3h4/rAaBNh8zjSXjTFYLBaQUmI+n0MIAeccoihCr9fDaDRCp9PhAIR9F7StGiIA0FqnrVbLZ1lGaZpSHMfh5ubGLZdLbIMPpGlKV1dXiKIofPPNN24+n/tf/OIXPmxetIGDEPZdcQDCGGOMMcbY0+js7Ez80z/9k/if//kfBSCqqiqNoqgtpewJIYYAJu12ezoYDE5ns9m9brd7EkXR0Dmn5IZK01RGUcQBCPtWDqs4AKCua6zXa8znc1xeXmK5WKCua3jvIaS4dV8QnoQhe4/XBCKHRwgzxhh7/xzO/TgMPvZv12ybzwnnHIqigHNud19rLVqtFsbjMbTW0FojiiJuhcW+l712WCqKIpJSOmNMVde1K4rCE5GvqirEceystbXWujo5ObGPHj1yn332mQfgt69p/mWGfWscgDDGGGOMMXbbrvIjz3P16aef6vV6ndR13Q4h9KIoGiZJkrVardPJZHJnMpnc6ff7WbfbHSZJ0tvO+yAiIiHErQGQjD2Lc27X6so6twk4iFBVFfI837W8KoriSaAB2oQeTbsrf3zOR6MZes4YY+z99rxZIMeu22+JZYyBtRbbodSw1sIYAyklut3urvojjmNuh8W+MymlEEJEUkoFwFlr6263WzrngveenHPBORestVYIURdFUdV1ba219uHDhw6A/d3vfuexq3tl7MU4AGGMMcYYY+wJOj8/JwA0n8+VUkp3Op3YWtvy3neqqhpEUTQej8ezyWTy0WAwuDsYDGadTmeQJEkriqLoTT8B9m6y1qIoCiyWS1RVBWctiAjGWpRliXy1Ql1VsNYiIGzCD2wqPgK2VSMBRwegNzj8YIyxD8u32e8f3sZ7v2ud2AQgZVlitVrhr3/96y4QGQ6HaLfbHICw70psq4ek1jpN07Q/GAyslFLEcSxvbm5CnuehLEsrhChDCOuiKAwR1dPp1PzhD38IX375Zfjyyy+Jq0DYt8UBCGOMMcYYY7eJy8tL+dOf/lQqpSJjTBpCaAshekKIQZIk2Wg0unP37t1Per3enU6nM47juKWU0m/6B2fvLmst8qLAxcUFlsslyrLcLSo551CWJay1mxsHwIfbcz32g4/9LfuWjoRF4daXn/TRZ4yx98Vhq6yGEALee0gpd5UhRVHswpCqqnatsOI4fhM/OnsPCCF0kiQdIYSKoiiO4zg2xviqqlwIobLW5gBy732tlCLnHKbTqX/w4EF49OhRAFeBsG+JAxDGGGOMMcYAnJ+fCwACgLp37552ziVFUXS01t26rsd1XU+MMZlzLiOiLE3TrN1uD9M07QkhJBGJF30PxvbttxZZLJe4ub7Gzc3NLgDR+kmmZo25dVTuYYXHsYoP9gxNmAEc7Yv/lCYM2RsifCto4lCEMfaO258T0lwWQtz6XGnmgwCbfWar1UIIAWVZAtiEJkKIXWsspXjJkT3fth1WLITQREQhBOr3+zUAr7X2AEwIwVxeXoKIcmttsf19u/rss88QQrBE5N/w02DvAN4bMcYYY4yxD14TfoxGI7ler7WUMs7zvE1EPWvtsK7rzFqb1XWdGWPG3vsBgK4QoqWU4kMf2fdircV6vcZqtcJiscDNzQ3yPEdZlqjrGs45CCGAEBAAhIPw41i1B4cgL7Bd5GuW+Qib1HM/wtgPRnaHlwqxOb9/PYcgjLH3xG6ft1ft1oQiQmyO72jmgjTtsK6urlDXNZIkQQgBSilEUYTBYIBOp7OrHmHsOQQRCSkloihqee9Dv9+vhRA+SRK/Xq+rPM/ruq6D9z4yxihrLUajEQaDwf5AdA5B2HNxAMIYY4wxxj50hG3bKwC7mR9E1DXGDEMI07quT4wxU+dcVlXVqCzLjjEmCiFw1Qf73owxWK1WuLi4wHw+x3K5RFWWt4aVb2Z7hFuVHw1ud/UdBYBIoGluJbZBiAAgiTbhyPbyLtTYVn+E7baZuhoA+L3gg0MQxti76liLv8PzTUVIoyxLPH78GNfX15BSwlqLKIrQ7XYBAFprpGn6mp4Bex8IIVQcx2mv18uiKJJFUcirqytbFIVdrVZERBEAGUWRr+vaL5dL9/XXX/sf/OAHNoQQeB4Iex4OQBhjjDHG2AdtO/RcjMdjHUVRTESpMaYdQujVdT0CkEkpp1EUTZVSk+FwOGy3212tdUREPPmTvZC1dndqQgwiQp7nWK1WmM/nWK1WKIpiN8ujaT0SDoaaPysEYc/RVH0QbcKPsA0/QkDT906EAAoBsqkOCc1/aBt6BHgSEAA8PQk//N6/J/9LMMbeRU3Asd8G69hny34AYq1FURS7+zYBiDEGrVYLWutdOyylFFeDsBfaVoJESZIIIYQXQjhr7doYU1tryRgjvfew1lpjjEvT1H7zzTf+66+/xuPHj/ePUWDsKfwHG2OMMcYY+5DRF198IQHoXq8XhxBaZVl2Qwg97/3YGDO11t5J0/S03++fTKfTbDabjSaTyWA4HLbSNI201vw7NXsm7z2MMSiKYlflkec51us15vM5FosFlssliqKAMWZzpyPtrZ4394MXlZ6N8KTSgwBQ2PwRLADIEDYn76FCgAoBwm+uEyFABDwJSEAQggDahCX71R682sIYe9c1ITHw7GC9CUCa220Xo1HXNYwxcM7tWjfuf15JKSGlvBWgMHaINoQQQgkhBBEpAEIIIZRSkoiC996WZWmUUk4pZQE4pVRYLpf+/v374eHDh2/6abC3FP+xxhhjjDHGPmTiZz/7mRqNRrFSKvXet621vRBCv67riXPuxFp7p9/vz6bT6fQHP/jB+M6dO4PpdNrpdDpRFEVS8F/07DmccyjLEjc3N/jLX/6Cy8tL3NzcYLVa7YKPsizhnLsdbuDpmR/A0/M+OPx4PrG3FSFAgjbbXfixCT6k95BN+OE8pPcg77fzQWgbomy3e3NZmsHojDH2vmg+V461xNrfNqHG/pwQYFMdUpYlrLVQSiFJEkRRxAEI+9a2gZxQSkVaax1FkfLem7quq/V6XQKwRGQBuDiOXa/Xc/fu3QuffvopHj58yB/K7CkcgDDGGGOMsQ8VnZ+fyyzLIiFE6pzrGGN63vtRCGEspZzGcTzrdDp3ptPpdDabje7evdsfjUbtXq+XNOEH8Qo0OxBCgHNutwi0XC5xfX2Ni4uLXehRVRXqut4NO38q2MDxqo/d1/eO1mW3NUPOxfb/kQQ21Rz+dvAhvYd0DtI6KGchzJMTWQvyHnD+SSWIwK32WCGE3WyQ3SyQN/OUGWPspaLnhLtN4LEffuxaAW7bYTUD06MoglKb7vtVVaEsy121CIDdYzB2oKkG0UQkAKAsy3K1WlXz+bzCpvLDAXAhBBfHsV0ul77f74f79+8ThyDsEAcgjDHGGGPsg7OZlUj02WefyTzPk/V63amqqh9CGDjnJt77LEmSk36/PxsOh6ez2Sw7OTkZnJycdHq9XpKmqebwgz1LCAHGGKzXa6xWK9zc3OD6+hrz+XwXfjStQprw49jJ783/2McvuyO2bal2Rydjs7AmtmGSwqbllQoB0jXBh4U0BtJaiMqA6hpU10BVAcYC1kLsqkDCkwoQIgQEBBACYVMFwjNAGGPvmd3spINKkP0qkMO2WM3nXzPzSikFIoK1FnmeI89zlGUJ7z2UUrsghbF923ZYUgihAZC1NuR5vp7P59VisaiFEA6A01o7KaVzztUhBF9VVciyLDx48OBNPwX2luEh6Iwxxhhj7IMSQqDf/va39Pnnn4vf//73KkmSaLlcdgAMQgiZ934mhDjpdDqns9ns9M6dO9PJZDLs9/udTqcTKaX4L3X2XN57VFWF6+trXF5e7oIPYwyIaLcg5L3fbQ8Dj2OVH+xpTbXMboEuBAjaBBXYDjXftL5qKj78JvAwFsJawNSgbcVHMAbBOQTnACFASgFRhBBpiDiGTJNN7KEUPBG8IPgAQGyOevbAJoQBD6dnjL1f9gelH17XhCJNJYjWGsCmFdb19TXKsoSUEt57eO/RbreRZRmEEFBK7SpEGDsmhCC891Fd1z1jzMR7v/beeyIK1tpARC6EUBpj3L179/z//d//4auvvsLZ2ZknIv4wZgA4AGGMMcYYYx+QEAI9ePBAfPbZZ/Lx48fSORdXVdXy3ncBDKSU4yRJpkmSzMbj8UmWZZPpdDoYjUbtNE1jrTXP/GBHNQGJkmcwAAAgAElEQVRGM/NjtVphPp/v5n3Udb0LPPb5gzkfh4PNeSH9QAgACESbdlOiORJ5+/9MgEAhbKo2Qti0v/IBKngIYyGNhbR2U+1R1Qh1BTIGqA2CqeGtg/ebAARSQiQJZJIguE04JbY/g5QKHoAXAiFsfg6xDUH4X4wx9j7ab4t12CKr+cxqWlo1n4fNnKumNZZzDp1OBwDQarUghID3HlprrgZhzyKISCulOlEUDdvt9hqA9d5b51ztvS9DCHkURfbq6gr9fr92zhEAG0LgEIQB4ACEMcYYY4x9IJrwA4BM01RdXFxEZVm26rruAugR0TCO43G32532er2T6XSaTSaT0Wg06nS73VQ3hzQydoT3HsYYlGWJPM9xc3OD+Xy+m/nhvT/aKuRZLa84+DgibAaS06bEAsCTAGQTQAACYRt8bLfboeZkLZSxkLV50uZqXQJVBV/XCFUFby2cMXDBbwIQrSGNQTAG0rnt9yJQAIQGCGo7G4TgQZDb4ei+GZDOGGPvmf3Pr6byYz8UaapAmlMz78MYsztvrYXW+lYA0ul0eFA6O4qIhJRSR1HU6Xa7xjln6rq2xpjaOVcS0dpauwoh2CiKsFqtxHA4rP71X/8Vq9XKAnxsAuMZIIwxxhhj7MNARERZlqnHjx9HZVnG3vu2975fVdXIGDOVUk57vd7so48+uvPRRx+dnpycTEajUbfT6SRKKcWVH+x5msqPm5sbXF5e4vLyEsu9yo/GfgVIU/1xeJ49jbZVFtuRGxBEkNsB5zIEKAA6ACoEKO+gnYe2HspuQg9V1aBiDSoKYHvyeQ5fFHB5DpvnMEUBU5YwZQlX1/DbHva7hb5mCjoJeCKQlCApABIIhN0ckP2h6Iwx9j46DD4Ov9Zs98/vX+e93w1EDyHshqXzsSbsmG27NBFFkYiiCACcMcbVdW2dc1ZKaaSUQSlFcRxDCBG01qEoinD//v3AQ9EZV4AwxhhjjLH33vn5OZ2enso//OEPmogSAGkIoeecG3jvJ977SQhhorUe93q98XQ6HQ8Gg36apqnWWhERhx/sKU3VhvceRVFguVw9mfuxWMBt233sBxvN+WNtr5rrecg5ngw1B7aVH9hrbdUMJd+0txK7VlceMoRNtYZ1EM6BnNvM+igrhPUaoSzh1yV8uTm5soTdVoE4a2GdhfUekBIURdDWQjkHbP9dFABBYlMNIgWC2AQxYVsdEgAEAleBMMbee89ridVUdgCAlPKp+6zXa1RVtQv/t4vWuzlZ3A6LNYQQpLVWnU4n1VoLrXUAYKy1ZtsGywohKgDCey8BSKUUoigKaZr6zz//3GNTBcI+YByAMMYYY4yx9x0BEFEUSaWUTpIktta2rbU9Y8yQiMbOubEQYiSEGMRx3G+32512u92OtoeZMXaM9x7WWlRVhTwvsFwuMV8ssFytUBTFreHchwNkn1Xt8UGHH/tHE+/Cj3ArACFgN99DYPMHLXkPHQKE9xDWbQOQzZBzMhaoa6AsN9UexfpJEFKWcFUFW20qPnbtWYBdABK2AVcIAUJKgAhKCEAQSElIpRC8hyQJT5ufze+FN1zVwxh7nx22xGrOH2uR1WhaYllrIYSA1hqdTmcXeLRaLW6HxXaISBCRiKJISSkFAF9vGACuqiqznQMCay2UUijL0tV17dbrtZVSuvPzc//ll18Gngfy4eIAhDHGGGOMvc/o7OxMAFDee01EcV3XLWNM13s/tNaOq6rKQghj7/3QGNOz1ibOORVC+IBXotm3sWl7VeH6+no38yPPczjrNgs3B9Uex87vX/ehhx/UhB7YBh7N9di2wArhyYyPEEBus5Xeb4acb8MPMgbSWIjtcHNU2+qPIgcV6//P3r30xpFe5wN/znnfquorm82rRM0YsBEEhhQgCJxNgAA2gqyyl/f5JFG+hj+ClQ8xWWSZ7DzLAA7imVgjkexL3d7b+S+qqtXiaP6xHXskdZ8f0GDzIopNUurueuqcB6hrxLpGaFv4tkFwrruEAJ8iQkoQY2GKApLS7msI1nZfozUw1oCyrLuOLrAR5q4YvV+FlYDu7RqCKKWOwMNS9P37tf0OrOEy9IVst1v85je/QdM0aJoG19fXmM/nsFYPWap39UFIfnJycmKMwWw2481mI6vVyrdtC++9MHMSkSAiYbFY+DzP4+PHj9PPf/7zYRJE75SPkP5vopRSSimlDhU9f/6cnz17ZgDYu7u7whgzjjHOYownKaWliFww84W19jzP86Ux5gTAmIgsgCM+Gq32Dauu9ovKAfSTHyVWqxVub2+x2WwQ+rVXTAzB2+mB7wo+BkcffgC7iRmSLuSACHhYd5X6CQ/0L+NwiTCpfxkjTAgg57uy87btCs/76Y9U15CqQmpqSNMitS2SaxGdQ/QeIXhEEUQRwFhIil3wQQQmQujXshhrgSzrAxDbLeNiRqIIw4xEjCQJ3L/UEEQpdSzed7+2H4IMwcd+ADJ0gYQQAACj0QjWWhhjYIfg+ZjvI9UOM5O1NptOp9Msy0xRFGSMiSGEVkSGgCMCcAAcM7d3d3dxuVzGZ8+eRQB4+fKlhiBHSAMQpZRSSil1sJ49e0YAbJ7nRQhhIiKzEMJCRJbe+wsAl1mWXc1ms4vJZHJ2fn5+MplMxtZaQ/psW/VSSnDOoWkahBCQUgIRwTmHzWaD+/s7rNcrVFUFYDhQ8/7n1kOAcvQTH3t2wQe6dVYEwKBfc9VPflDsOj04JVAMYB/Avn9bCDAxgLzvPs57oG5ArQNXFaipQXWN2DRA6yBtC3H9S++AECDeQ2LoV24JxFoQBEIMMdxNd2QZkjFI1iBZC7YZyFiYvhA9EXUTIMYgESOKgIm6lVjQoy1KqcO3f7823M89XIclIrDWYlhZ5L1HXdcQEWRZhvF4vCtKH9Zh6TSI6pExxjKzNcZkzEwppeScC8YYVFUlTdNE733rnPPM7LIsi/P5PDx9+tQ9fvxYnj17Ji9evAD0bvmomP/9Q5RSSimllPr0PH/+3Pz4xz+2eZ6PRGRKRLOU0mkI4TyEcBFCeMTM17PZ7Pr6+vr8yZMny5ubm/nl5eVoPp/nWZYZZtYj1ArOOWy3XcH53d0dVqsVNpsNNps1ttstttstutULAcC7xeb7gcfw8tjDD+knPoaeDOonLBjdE1QLwIjACmBTQi4CGwKyEGFcC9u2ME0Lruou4KgqoCxBdQVsS8i2BDYb0HoFc3sLc3cHur9Dqmr4toF4j+QcxHkghi4ACQEkaReAMAiGGWwYhhiGuwszw7CBNRbMpiv37TtLQH1Qwt1ECNAdXTniH7VS6oi9r//j4VTIcH2/9DzGuDvZIMsyGGOQZdn394Wrj1n/sIFob50aGWNMlmVsjJG2bX0IwYUQfFEUfjQaxfl8HheLRVosFvLrX/9afvazn+GLL77QAOSIaISqlFJKKaUO0nK55LZtbZZlhbV2EkKYxxgXKaVlSumciM6zLDufzWZn19fXpzc3N/Pz8/PJdDrNi6LQ8OPI7QcYw6qr169fY7vdomkaGGN273d9f8Tw5/b//PvWXh1r+DEEH7uej/57MUx7GKALQmJChm7qw6TUlZr7AGod4Fpw6yB1DWoaSNt2JefeI4UAeA/yHqj7cGS9ApdbkHMgNmBju4AjpW5dVoxADKCUECX1PSPoVlf1fSJsLdBPjCDLINYi2QwmsxBruoN3xnS9IdYgG55mD10g/e2W7pugiYhS6mjsT4AM05MPe0GMMbt1kU3T4PXr12jbFs45FEUBa+0uCNF1WGoPM3M+Go1mzGz6qSJ3f39fxhi3IYQmpdTEGEPbtp6IEoD09OnTYQXWd4/rqoOjAYhSSimllDok9OLFC/rVr35FP/7xjy2Awns/EZGZc+4kxrhk5vPRaHRRFMX5bDY7u7y8XJ6fn8/Pz88ni8WiGCY/9An2cYsxwnu/t+bqHuv1eheADOs4iAgxRsQYMUx/AN/u+TjqyY+99SfdhAXA6IcmksBQt+bKAH2huYBDhE0JJnQrrqh1INcCTQv0Ex/YbrsQZAigUtoFIFTXoKoEb9agsgTFCJtlyGwGECOJIMWIlBJijEgpIojAo1scnoiQYuxCmNAXqjdNv96KAJt1a7DYQPoVWGwt2BoYayGmW++SIO8eXTnGn79S6qjtBx7fFYIMAUlKqV8n2b3v5OQExhgwM/I8R5ZlOg2iAOwmhwwzF0RkYoyeiLYA7kMIqxhjFWNsYozBOecARCJKP/rRjxIAEREhIg1AjoSuwFJKKaWUUoeCnj9/zn/5l39pxuOxHY1GI+/9NKW0dM6dee8vvPfXWZY9ns1mj548efLoyZMnl0+ePDm7uLiYLBaLvCgKa4wZ0g89UnnEmqZBWZa4vb3F7e0t7u7udquuYn/gHMC3Ss6/a+rjGMOP3cTHsOoKgCGCkX7VlQgyADYJspiQxdhdnO8ujUPWtrBtA1PVoLICbbtQw9zeIXv9DfjuDrRaITUNUHddH3a7Qb7dIC+3MGUJ4xw4BEASqJ8oyYJHFj3yEJCniCIl2H4ChKSfRCGCIQITg4HdZbgtzNwFGtwFIDAGnGUgY0DGQNCdWtr9HpCeZqqUOnoPV189XIn18D506AkJIbwTgiiFt6uwGAA552JVVe7169d+u90G51xi5iTdL1RMKYU8z1NKKb1+/Vo2m43c3Nzgiy+++NC3Q30PNABRSimllFKHgH75y1/yzc0Nl2Vpr66uMhGZpJRmKaWzEMJFSumSiK4mk8mjs7Ozq88///zqyZMn59fX1/P5fJ7neb4ffqgjNay1qqoKq9UKr169wt3dHTabDdq2fafMdb/Q9X2X/fcf46/VLvzYW3XFSWCku2QAMnkQfnjfXVrXd3004LqGqSpQWYLLErzquj2y16/Aq3vwdoMUAqRtYdoW+XaLvCqR1RWM811xeh9umJSQpYgsBuT99UIS8pRg+vVXuyJ7YjD1YcdwkE7eXkefk5JhkLWgLOumQPKsW4mFbv3VLvig7pNpEKKUOmYP11gNHSCD4fqwgnIIQIqiwGg0eicAOcb7VvVtIiJt24btduvv7+9DXdchxpj6CY8kIiGl5FNK0RgTmTkZY+Szzz6TH/7wh9oHcgR0BZZSSimllPrU0fPnz/nu7m4XfpRlmaeUxk3TzEIICyJaTiaT8/F4fHl6enp5eXl5cXFxsVgul9P5fD4yxrCuvVIhBHjv4b3HZrPBarXCer3ehR8Pfz/eV3S+f/bqw1UfR6G/7bvb3H8Phm4NlrcBiI3duisTAmyM3bor72C8h2kd4BzYeaBtgboCVzVSuQWt1zB3t7Cre0jTIIYAM3IgZpAIbNvAti1sDN36reFrSgmG9gKJB1e4H/oSJHAiMEWESEgUAP92giMCADGiMQAbILOgPIcdjWDGY1CIiDYiGYMg/TqtvlwdBBDo4WIspZQ6Gg+L0Ye3DUHIcL8aY0Rd17uPmU6nu/BD12GpB4iZTZ7no9lsduK9b7Is8ymlAMCHEGprbUVEDoAriiKmlFJd1+mnP/0pdB3W4dMJEKWUUkop9UkTEfryyy95u93a6XSa13VdABjXdT0HsKjr+no8Hl+dnJxcP3r06Obx48ePrq6uLs7Pz0/m8/l4NBrluvZKiQiccyjLEvf397i7u8P9/T02mw2cc4gxvhNm7IccD4OPwbEFH92qK9r9I2L0q6SGfg8BrCSYmGBjQpYSrO/WUFnnukvbwNZtN/VRN6CqAlUVsN6AViuY1X1/WcGWJahtQKELOjhG2OCROQcbAzjGXfgB9BMpfSBCIiAMl/4fPr1db0V9UDFUpO4meYabC4FQtwKLbN//kecwef52AoQIsY86EgAZ/os5pt8LpZR64He5bxzub4cTDIB3TzJgZlhrYa09rvta9V1keDwGgLMsE2MMUkopdlprbcvM3hgTAETvvZyfn8ff/OY38i//8i+iUyCHTSdAlFJKKaXUp46ePn3KX375pd1ut1lRFKOU0oSZZ977EwCLLMvOZrPZ5c3NzdWjR48uF4vF+Wg0yvM8z/SJswK6IGOY/Pjtb3+L+/t7VFUF7z1EBMa8PXfs4aqr4Un3sPLqmOz3fAxI+gChn/qgPgDhYeIjxm76o5/8sM7DOAfrPahpu86OpoE0DdC0iHUN3m6A9Qp8fwdTlV2xuXOg1IUcuWu7v1QEnBJ476DZ74oBZJB+VdbbiRBg6PLoB1z6tVZiDMQwqMhhRiNIXYNcCxsCUkwwlGANIfbfB9Ovddn1gnTVIEopdXSG+8uHJxU8XC85vL9tW9ze3sJ7v5sKyfMco9FIAxAFAJRlmZ3NZuMsy+x0Ok339/cSQoje+zaltIkxrq21tfe+McY4Y0wIIfjLy8v09OlT/SU6cBqAKKWUUkqpTxn94he/MOv1OsvzvEgpTURkHmM8aZrm3Ht/0fd/nBljlrPZbHFycjI/OTmZMDMbY/QJzxETEcQYEUJA27ZYr9e4v7/HarXaTX4MfpfJj2Hl1dF4UHKOIfAAwNL3ZaQE0wcS3K+5MiHAhAjyDuQD4Lp1V6l1YOcQmwbStEBTg5oGqCrwdgvarMHrNbipQG27W28lADjG3VIp2pvU+H3svvb+c0AiJPUTIUngjSBAsPubmAFjEKsKsSggkwlQN6BxC2MzWAAZDCIzhIf1Wv30CET7QJRSR+194cd+z9Z+GXpKCXVdI6WElNIu+HDO7T5+KEkf1mMd1f3xket//lwUhbXWGiKaiUhq2zZmWebKsqxFpDLGOCJydV2HPM+Tcy4CSHd3dxH9hkt1mDQAUUoppZRSnyp68eIFff311wZABqAYj8eTGONJjPEshHARQrgMIZzFGJciMieiaZZlRZ7nujRaQUQQQkBVVViv17vLMPkRY4Qx5p2DMMPL9629OqqDLdKNeQxrpbifvjAgsAAMeRt6xAhyHhQCjPdg77vXnYM4h9S2QOsg3nfXmxbUNDBtA6prcFUB5aYrQa+rLjiJb49TDOHL//m7L2/XYRkCMgESUre/qg8r0nAhAoxBaltI20KaBqmuuymQpukK0Ym6qZKsX7Y1/H4IkLQHRCmlALz/vvN905TDpGZZlri7u0NKCdvtdvexo9EI8/kcp6enuxVZ6mgQd1OWhpkxGo1GMcZ0dnaWiqLwo9Gorut6671vmqZx1lovIkFEvLU2fP755x67pZfqEGkHiFJKKaWU+iS9ePGC0Z2snU+n0xEzT0IIp9778xjjdYzxOoRw7b2/KorifDabLa+urk4Wi8VkPB7nH/rrVx9ejBFt2+L+/h6vXr3CmzdvdpMf6cEKpf8t/Dgq+6tK0PV8kAgsUd/zIbAiyGJCFiNM08K0LUzTdL0eZbfCCmUJ2WyRNhuk7RZhu0XcbBHKEqmqkDYb0GYNu1nBlluYpgZ5D0pp9zX8qQy3zfRhDqE7NXQIQLot4wwwd/0fxiArCmRZBmMtyFiAqVuT1X8c+imQhP73CHqkRSmlBvsrr96nP8C9C0KqqsLd3R3evHmDu7s7VFUFZsZkMkFRFO+srlTHhYhgjOE8z7OiKMham0IIwXsf27aNzOyJKBBR6IOQ8Gd/9mfhiy+++NBfuvoT0f8NlFJKKaXUJ+fFixf81VdfmSdPnmRt206Yeeq9P0kpncUYL0MI10R0Za29nk6nF8vlcnl+fr64urqaLhaL0Xg81tMCj9T+2qu6rrHZbHB/f483b95gu92ibdtvTXXshx1HGXwMK0mkO4Y/TEmwdE8oTeo6M7K+3yNLCTZGZCHAtG4XfJi6m+gYis2lLIGqRNqWSFWNVJWQupukiFUF1BVMXcHWJUzTgMP3E34Ae+EO3tZ0DEXmXXV6X2rODLIWxlrYLIPNMhjbhSDC/G74QdT/+bchivSTNEopdeze6ZJ6cH24AG/vx9u2RV3XKMsSdV0jxghmRlEU73w8Mx/XhKbarcQyxlhjjBBRAhBFRJg5MbMDEGKMPsYYRCQYY9I//MM/0F//9V9DC9EPjwYgSimllFLqk3N5eckXFxcZERXz+XzqvT8homVK6cJ7/yil9DjP80fT6fTy8vLy4vr6+vT6+np+cXExns/nWZ7n+jj4SIkInHOoqgqr1Qp3d3dYrVZYr9domgYxxm+FHO+b/jgmNJSLg0DoXhoQjAiMACalt6FHH3zk3sP2ZeamqmDqGrw3+YHtFtJPgEg/8SF1jVjXkL4AnZsGpq6RtQ1s8OAYv5fwY3e7hwt9u6s8ARAmCDHYGLAxXe+HtbDGgJhBbABrQNy93gUgXXAS9z6HHpZTSqnO/hTIfogxvD58TIwRzjl479G27W5yc/iYYYrTWgtjzG56RB0HIqI+ADHMPLzKxhjKsgwpJRdj9E3TeGaOo9EofP7555GI8JOf/ER+8YtfHNcDvSOgZ74ppZRSSqlPznK55EePHtmiKIqqqqYichJCOA0hLPv+j/PJZHI2n8/PfvCDHyyvr6/nZ2dnk5OTE6vhx3FLKcE5h7u7e9ze3mKz2aCqSnjvdwdeHoYfw+XhWqxjsJv2YO7KxYVg0BeNi3QhSIiwKcHECA6hLzkPYO+BpgHKCmgaSF0Ddd1dr/qXTYPYNECIkBAg3oNiBHmP5B1SCMAH/r4zAAvBuC91J3ThRYwMiQHwXYm79LcxFQU4y0CZBecZYA2kT1ISAZEZLALmvUmSlHQdllLq6O0Xoe+/bf96v94IAN45aSHGiNVqtVuP5b1HlmXIskz7QI4YM2dFUcyIiLMs46IokFLaeO+rEEIFwDGzq6oqzmaz+j//8z/ll7/8Zfr5z3++23ipPn365E8ppZRSSn1SRIT+4z/+I2PmMYDZXvBxzsxXeZ5fTyaT6/Pz84vLy8vlD37wg5PLy8vJcrkcFUVhrbVEugvhqAzhhfceTdNgs9ng7u4O9/f32Gw2aJr2vZMfKaWjm/YAsFt5xXhbcN6tvOonPvqOj7cTHxHWOVjvkTkH27TgpgFXNbiuQWXVhSDDBMh2C6rKLiyoKqBtQa67cOtA3sF4DxMC8hiQpwQj6YNNSuyvw+reAHgiRGIkZhhrwYZh+wkQYwzYWpAx4Mx2EyCGAWIkIiQiRGakYbxkn67EUkodufeFIMPb96dC9ldcDfff3nt475FSgjEGeZ6/0wXycKpEHYVhGiTrf7diWZbbsiybuq5bZg7MHIwxcTwex+l0Gi8vL+Pf//3f4+XLlx/6a1d/JBqBKqWUUkqpT8rLly8ZgDXGFDHGSYxxnlJaxBiXRVEsZ7PZ2Ww2W56fn59eXV2dLJfLyWKxKKbTafahv3b1YaSUdp0fVVVhvV5js1lju92irmukFN/5+IedHw/fdtCGvg8M65+6gnNGF3ywCKwAJkaYGGFD7MIK78Heg50Dty3IOaBpgabtQo6+9wNlCa5LpKZF9B4UAsQHmBhAPnTTHymBU4JNESZ1r3/w7wm6swctAVbQTbykhBgjKESQDxDXIjUNUp5D8hzIM1BTgKwFjIEQwzCBiWCYYYiQ0K/Xoq4jRCdBlFIK/9+Qou93eOc+2VqLEAJCCPDeg4iQ5zlGoxFEBKenp5jNZhiNRroO68gQERNRzsx5SskZY05SSqcxxqVzbsPMLYBGRFyM0TOz32w2/vLyUt4XxKlPkwYgSimllFLqU0EvXrygu7s7XiwWtmmakYjMmHnhvT9LKZ1PJpOL6+vr8ydPnpydn58vFovF7PT0NM+yTCefj1hKCU3T7KY+7u/v+/UYDiIJKQm6mgvZffz+KqxjCT+ov43UH/Afrhugm/yAgFNClgQcAmwIsD50XR9tu7ugaUBtH340DaiqgaoCyi3sZt11gHgPEUBS/zmDRx6HwKNbr8WSYJBgIB9NT8ZuJRj6SZgk4BhBIQDOdyu9rAUbA7IWnBfdJAgTDAGGCdZwtzoMhMQMSgkJQBLR8EMppb7D++6Hh3VY+9MgIQSklLBareCcw3a7xdXVFW5ubmCM0XVYR0xETIwxd87NvfenIYTSe++zLGvzPPchBFfXtSuKwtV1LS9fvhT0lV0f+mtX/zf6RFAppZRSSn30RISIyDx9+tS8evUqb5pmFkI4jTGeE9H1aDS66tdeXT9+/Pjq5ubm/OLiYn56ejrWtVfHY3/VVVeO2hWk1nWNsix3Ach2u0Xbtggh9AdU5L1hx1EEH8PEx97aK8aDdVcxwUqCGQKPEGCdh2la2KaBrSqYsoQtS/BmA7vdgrZbYLsBlSVkW4KqErzdIttsYKoS3DZIMUJiN/VRxIAiBeQpIpMEi27NlkE3ffKx/ONNREjoS8ypKzY31PWiGCJY9EEREdhYkLUgwxBiCDPEGIgxiNb0b6PD/x1TSqk/gu9aizW8ff8iIgghoG1bpJTAzCiKYleI/nCNljoOMcbgnItlWbbe+wAgWmuTMSYQkffee2ut9957ZpZf//rX+Md//EfRVVifPg1AlFJKKaXUx4xevHjB//qv/2rOzs5MXde5tXZU1/UcwNJ7fzkejx/NZrNHy+Xy8dXV1dX19fXl9fX1YrFYTCaTSWGMYQ0/jkOMEd57lGWJqqpQVSWapkVVVbsAZL1eo6qq3Rmi+yHHfsn5sRyUpn4VyLurrgBOfc9HSrAxwvg+/PAetmlhmgambmCqGrzdwGw2MPf3MKsVzHoN2mzA2y243IL67g8uyy4saRuwc0giQBKYlJCnuAs/jKRu3dZHFn4AXWG5gLrichoK0vuLoAuKUoIBgZhB1kKYAO5WXIm1SMZA8gzCDHB3CwXd9IfoFIhSSr3X8FBuPwh52AsyvG0IQJqmAdBNhlhrwcy7AISZ3+kHUYcvpZRCCOKciwCknyBKIhJijIGIWgBuMpm4PM9lsVhI27by/Plz9NMg6hOlc19KKaWUUupjRl999ZX5m7/5G5NSyohoVFXVxFp7UpblMoRwNh6PLx49enR5dXX16Pz8/PLs7GwxnU4La60+qz0yIQRUVYVvXr/CdrNF0z2XjOUAACAASURBVDQwxvQHQuJu8mO/3HwIQIbL/uqrQ0d4u+5qKDvf9XwAMCmBvYfxAcZ7kHPgtl935RxQNxDXQjZrYLMBr1bgquzWYIUACQESIzhGoF8RZZwD9YXzeYow1IVONnV/78cUdrwPo5vwKKT7/iQIEASQBIoB7Lsyd4SIBEHM+gCk7/iQLANZCxNGyIztQo/+koDdFE46kt9BpZT6Qzzs6RpCkKHfYz/YSClhs9ngq6++Qtu2cM7h+voaxhhkmdbDHRNjjBmNRsX5+flpURQ0nU7NarWSu7s7X9e1M8ZUxpiGiNrJZEIiQovFAp999hmkG0f/wKVk6g+lAYhSSimllPpY0fPnz+nm5sZsNps8y7JR0zSzlNI8pXSWUjoLIZwbY4buj4uzs7PlbDabZ1lmmVkDkCMwrL0awo/1eoU3r99gtV6hrmswMZjN7mzQYe3VwxBk//MdOtp7ydL1bRgicBJwirBJYEOACQHGeZih36NpwVUFKkugabqSc9eCNhtgvQLd38HUNahtgCQQSUA/5dG97MrN0U/aUEqww972TyD8ALArQ6d+RZck6m5bjCAmkGOIc5CYEJgQ8ryfGummbSTPwXmBLA7l7t3vZhKAZW/RuEgXmiillHrH+05U2J8K4b3JxkHTNPDew3uPlBKyLNu9P8uy3WSIOmxEZLIsK+bzOed5zlmWmRhjatvW9wXoVZZltbW2aZqGsiyjPM+lrmv54osvUh+CHP4DxQOkAYhSSimllPoovXjxgh4/fswhBFvXde6cG4cQ5imlU+/9EsBSRJZEdGqtXUwmk5PpdDobj8fjD/21q+9PjBHOOzRNg/VmjdVqhdVqhfV6jbqu+3LUbx/Y2J/6ePj6IW9MIwDopz1IhrJxAaXUdX7ECBsjsv3wo2nBdd2tsdpswOt1V2retkiuBZclzGYDXt2Dmhrs/e/0tZj+a/mk9GvCeO/1nTi8DAgiXRF6lndBBjMky4DRCDzxoBCBGCHRIFIXfKRhvZak/gAfPq79X0op9ZF4Xwjyvl4PY8zuJIm2bQF0gcdkMtl9jul0ijzPNQA5AtzrywFZRLht2+Cca0XEAVjHGMumaaqiKISZU1mWqWma5L2P//zP/6yF6J8oDUCUUkoppdTHiABwWZa2bduMmUcxxmlKaRFjPAshnDvnzkMIp865eQhhHGO0KSV99npkfPDYbDa4u7vF6v5+F3ykFMFmCD7e7g3vCs+/PfWxv0bj0Miw5mo4OxbdxAX3XR8cIzilXfhhvAf7AGod2LWgugZXNWi9hr27g7l9A2w2IOe6EvPWwbQNqG2BqNshIAIOAaaqIERgJEQmpKIAprNulZgPsHlCihGWGXGv74RBkC6p0hBEKaW+w8MQZP/6EGYMb7PW7l7fbrf4+uuv0TQN6rrGo0ePcHJyouuwjowxhouiKE5PTxdZlvn5fB6rqlpvt9uyaZqqrmthZkHXFRJjjP7p06fhQ3/d6g+jawGUUkoppdTHhl68eEEADDPnTdOMRWQaQlg45y5E5DKldEVEV8aYy/Pz8/Ozs7PF5eXlbDqd5nme60k+B25YYRVjRFVXWK1W+OabV7hfrbDebOBci9RPcnQrsAhD00IXduBb0x8HS94tEh/WXpm+w8KkBBsibOiDj7aFda4rOK9rcFmBqwq8WcOsVrC3b2BevYJd3cNst+C6gm2abkVWCGDRAAQAIN2KL5NSNwFiLVIxAkZjUDGCKQrAGJAxiBBIPwUyrMvqfiVJww+llPr/eN/Ux/s+Zr8oPaW0W4klIiiKAlmWwVq7mwI9xJMh1LcQEbG11mZZRtZahBDqtm3bqqralJKISCKiwMwBgHfOpWfPnskXX3xxwA8cD5M+OVRKKaWUUh8jBmBjjDmAUYxx6pxbiMg5EV1nWfaoKIqr0Wh0cXFxsZjP55M8zzPW/QVHIcYI5xyapsZms8H9/T1WqxW2223X+8H8ThnqEHCk9O66q/33HaT9Xo3+ugHBgsApgmOCDaErOg8B1LYw/YVbB25amKoCbTfgzQZmdQ9zdwt7fweuK1DQEyG/C0kChQRJEWwMeDIFmgbSNKCm6b7HWQZkFpk1iEKwTIhEXUhFhASByBDeKaWUep/9sOJhcLHfB0JESCnBe48QAlLfRzWdTnfvm0wmu0BEHTZmJma2xhjLzFFEvDHmIsa4CSGUKSVh5sjMPqXkYoz1Z5995i8vL7UL5BOkAYhSSimllPqY0PPnzxmAHY1GWdM0BYCJ934mIgvv/YUx5no2mz26vLy8vL6+Pr++vl5cXl5Ox+NxZozRAOQIeO/64OMW6/Ua96sVnHMQEVhj3imPHgYS3tf5ccgI6L4Pe+uvusmPrvPDptSVnHsPdg6mdaC6AtcNuO7WWUlVAWUJXq9g1yvYzRq82YBcC8T46fV3fF/2vy8CICVICBDngLYFtS2oaUFZBrYWLBmMNWBiGAxdIN2fFV2DpZRSv5P98GP/Pn44IeLhZIeIoK5r/Pa3v0XbtqjrGpeXlzg9PdUA5Dj0D5UIImJFpPDenzjnzmOMpYhEIvIxxpaZ68lksmVmV9d1AjBMh+gDoU+EBiBKKaWUUuqj8uzZMwJgU0q5MWbsnJumlE4ALK2159baq+l0enVxcXHx+eefn15eXk7n83lRFIW11moAcqCG8CKliLpusNms8c0332C9WaOqqm7lEBGstUgikPT+kvPh+iEjvLvyagg/SACOEUYExgcYH2Bb162vqmtQVYGrGigroGlAdQ2sVzCru276oyzBbQsKAXTg38M/FkJXNI/gQc714UcD1BUoy2CyDEwCQzkMEQz3hehMu1UsOgGilFK/n4eTIPtrsIaLiKBtW9ze3qJtWzjnYK1FnucoiuKd4EQdPBaRXETmRHQGoCEiLyJtCKE2xpQA1tba9smTJ/HLL7+UX/3qV9AQ5NOhAYhSSimllPpoDNMfV1dXWV3Xo6ZppiIyZ+ZFnuenRVGcTSaT88vLy7Pz8/PT8/Pz2enp6Wg0GlkiIt2AdbhijPDeo21brNb3uF91a6/KquwOWhgLYgb6FUIg7NZbpJSOI/yQbuiD+vEBA9p1fiBJ1/kRI7KYYJzr11w1XfhR18C27MKPqoK0LVJVgTZrYL0Bb7fgptbw4w8RI8h5UFmCyi2oKMCTCSTPQUUONt1BNsuMJNJNgBAhEQEpgQR9KbpSSqnfxXBf/77wYnisGGNEjBFlWe5WYo3HY+R5DiLCaDTSdVhHgoiYiLI8z2eTycR571vnXB1CqFJKZQhhIyLTsixdlmUpz3N5/vx5Vy6nZyl8ErQEXSmllFJKfTT+9m//1s7n8zylNPPeL0TkzHt/boy5PD09fXRzc/PZZ5999vjx48fn19fXs+VyORqPx9Zaa6h7lquHCQ9QSglt22K9XuH169d4/c1r3N3dYbvdwLUOSRKIuZ98IEiSXeiRHkyCHKpu0qMLP4auDwN0Zef9yisbAqzzXc9H3cDWNbgsu+BjuwE2G6T1BqksIVUFqUpwWcFWJbKmgfEOlLTk/PdDfShHoJTARDDGgLIcyCzEWggzEhNgDMQYgOltGTr0yIpSSv2+vqsc/X1vjzEC6EKTGCNCCAghgJmRZRmyLNMpkCPQTwaxtZaNMUJEoW1b75xzfT+IN8bEPM9TCEFevXolX3/9tdzc3EBL0T9+OgGilFJKKaU+FlQUBTdNkxVFMQEwDyGcisgSwNl4PF5eX1+f3tzcnCwWi+l0Oh2Nx2PDzPqs9ICllBBjRNPUWK/XePXqFe7v71HVFULwXfgB7kIPIhAlpDQEH93nGAKQgzyA0d8uItpNfjC6qQ8GYFICxwibEth5mNbtJj6oqoGqn/ioKqRt2b3eNBDXgpu2mwTxHqk/QKR+XwIKAdzUsMFDDAN5DsznkMkYaTQCrAEbA5NFmJSQmJAE3c+RgLQX3ukRFqWU+t0M9/n70yD706DUB9LGmN06rDdv3sA5h6ZpwMy7dVjGmG91iKjDwcyUZZmdz+ejLMvEWutEZLPZbDYxxk1KaRtC2DKzSynFPM/j3d1dtNamp0+fpq4TXVdhfcw0AFFKKaWUUh8avXjxgp4+fUpffvllBqDw3k9F5CTGeJpSWgJYGmMW4/F4dnJyMlksFqM8zzNjjK69OlDDmZjDgYj71Qr3qxVWqxU22w289+8cjOgOZghServy6qAnP/aCDwCgvuy86/ro1l2xCEyM3SVEcNvCNA2orICqhpTdyiupKkhdQYa3tS3YObB3oKaGCaGb/DjQb+WfGkmCCR4cI2JdIZZlN2UznULGEyDLwZmFeAtjbb/+imEgiAQwEeIQ4A2/03oQTimlfifvPk54OwFCRIgxgpmRUkJKCXVd7x47TCYT5HkOZt6tw7LWaghygPo1uibPcyIi8d5PrLUzAPMY4yLGWBZFsW3b1oUQQl3XPqUUAUQA6eXLl+ivq4+UBiBKKaWUUupD4ufPn9Pjx4/5yy+/NADyoihGMcZpCGEhIsuU0jKldBpjXIjI1BhTZFlmsizT5OOAiQi899hut7i/7zo/3k5+dLu6jelaLoYDGV3wsV+Y/nZd06EdsOgmPrpEgvvrLOjWLPVdHyYlGO9hQoDxEdQ0oKoCyr2uj7KE1DWkqpHqCqhrcNPCeIfMOeTBwXgPlgRNQP4Ab8eQQEggHwDnkJoGqa4hdQ3KMyAz4CyDzTKIMbApIdAwBdKvwxo+13AW84H9Tiul1J/SfhDCzLuXxpjd2wHAOYeqqvDmzZvd62dnZ1gsFu98vDoo1D+WNMxsmTmPMU6cc3Pn3KmI1N77sq5rXxSFs9Y2AFzbtmE8HqevvvpKtBD946YBiFJKKaWU+lDoZz/7GT979ozLsjTj8diGEAoRmcQY5ymlRQhhGWNcppROnXMnMcaxiFho18fBG3o/VqsV/ud//ger1QpVVcGHAIBg2ICJ3/l4gN6Z+hjWXRza+quh7IaIwP11FukuKYFCgAkB7D2MD2DngNaBmgZSlqCyhJRVdxlWXtU10DSgpgG3DXLvUDiHPHqYFLvP+2Fv9kEQSUjBI7ZNHzhV4DwHZxkkd0CWIRmDxAzDBMPcr3YjxJR267D0CItSSv1+5OHkZH99CEP2T6ZwzuH169eoqgpVVUFEUBQFRqPRB74V6k9NRCjGaJ1zI+fczDm3EJGmbdvaGONSSk2WZRWAhpm9MSb83d/9XXz58iVrCPLx0gBEKaWUUkp9CPT8+XN+9uwZA7DOuWwymeRN00ycczMRWYjIcjwen52cnJxPp9Ozy8vLk+l0OtorPFcHbFiB1TQNttstyrKE9747Y5P6Yml6N/DYn/jYX4F1SL8uBLxdf9V/L4bwg0J8G3w4D2pboGmAtgW1DqmqQFWFtN2C6qZbedV0wQeaFtw0MK6B7Sc/8hCQpbhbr6X+CJJAQkByDrFpgboGFQWQZ6A8A9ms6wMxBoYMLAgJQAIAZkCkW4cFDUGUUur3sd8Bsh+CMPMu+ACwW4lV1zW89wCA0WiEPM+RUsJkMtF1WAeMiMgYYyaTyWixWMxFxHvvvTGmDSE4Zm6IaJvnec3MfjQahf/+7/9OP/rRj4ZRWb17/ghpAKKUUkoppT6Ib775hk5OToy11hZFkTFzEUKYxBhnbdue9J0fy+VyuTw7Ozu9uLg4WSwW4zzPrQYgx2FYYxVj3O3n7g5UPPy4dwOPfQf1q9KvPWIiEABDBIOu/4Njt/aKfVd0Tm0LruvuAHvdIFXdeqtUlkC/eglNF5BQ24LaFtY5ZK5FHj2yGLrJj+6b+6Fv+cEQSZAYEdoWqW2ApgbXBUyeA3kOyguwtzB5DguDCMAyIwy/2xp+KKXUH+x9RejD2/d7QYbHE845bLdb3N7egpnhnMNyucRyuQQRwVo9rHpomBl5ntv5fD46Pz9PeZ7HsixD27at975JKW2Z+V5EtszcZFnmptNpOD09DQC0EP0jpf9SlVJKKaXUB/Hnf/7nFGPkPM+z0WhUpJTG1tqpc24O4ISZTyeTyenNzc3pzc3N6dnZ2Xw+n49Go5Fl5gM6qq2+y3BwoSgKNE3zTrghkvqXeG/wcZD64APouyHwdvWVhewCEG5boJ/2kLLsuj62XddHqqou/GhbkPOAa8Gtgw0BmWsw8h55CjCp+7zqj0wEEiOSdwhNA24axLybAjF5DhoV4DyDBA+TWRgCEjMkJQiwW9WC4XJIAZ9SSn0PHp4Y8b4QZHhbjBHee7x582Y3kRpC2E2EqMPDzFQUhVkul6OiKHiz2eD29ja9evXKee9r7/3GWnsbY1zneV5575vNZuOZ2f/7v/97/MlPfpL+979Ffd80AFFKKaWUUt+758+f81/8xV9wjDHLsizfbrdjEZkbY07H4/HZaDQ6H4/HZ+fn58urq6uTi4uL6WKxGBVFkRljWCdADtOw9irGiLZtUdc1nHO7yY/h4O/Q99GVnr9/8uPg9OuuCG+DD0oCA4GJCew82DmYtlurhLoG+sLzuN1CyrIv3W4gTQNyDnAO7D1sCLDeIw8BeYqwKXWf/0Pf5kO0C0A8xDkk5wDvIG0L6SdxKM/BeQ6TR9hkIEkA9EXoEKThZ9OXoyullPrj2O8EMcbsHnM0TYMQApgZi8UC3vt31m6qgzKswKIsy8ham0TEt23bMnPtnNsQ0VJEts65JqXkx+NxTCn5zWYTX758mQDED30j1Ls0AFFKKaWUUt+7Z8+e0X/913/Z6+vrvKqqcUppzsynRVFcnJycXE0mk6uTk5Or5XJ5fnl5ebJYLMaTySQ3xpgP/bWrPx0RgfceZVliu93uuj9CCA+mP+Sdl8dgd4YquvDDCGBEwDHChgh2HtS0oKqGDBMf5RZps0EqS8SygjQ1pGmA1sF4D/YeWR98FDEgjxE2RRjRgzp/KiICSRHJB0TXFdOnYgTOG0hRgFoHLhzIe4j3gM3Apl97JQIBkKjrBZHuE37Q26OUUp+qYR3WbrIOb+9rmRnA21Wc3vvdyRlD+KHn4hymvgOEjDHMzExEEmNMIYQ0Go180zRl0zRr51wpIq2IhKZpYkrJr9frCOyqu/QO+iOiAYhSSimllPq+0Zs3b8xkMrFt2xZ1XU/zPJ+nlM4mk8nFZDK5/uyzzx6dnZ1d9wXo474jRJ9pHrjh4ML9/T3evHmDzWaDuq7Rti1CCO+cbTkcfDj0EIT2Xg5rrwy68MPGiCxEsHPg1kHqBqmqIWUFqUrEsoRUFVLT9JcWaNtuTVY/9TEKfhd+mCTQmYI/MRFISkAMQAgQ7xGbBlwU3eqytgXaHFwUsHkGZB5kGNKHHon2ApB+BZakpKuwlFLqD/DwccQwUToEIMwMa+2uL8QYA2PMO6GJOlxERNZaO5/Px8YYzGYzv9lsytvb27WIbOq6blNK3lrrAbRFUbiTkxP/4sUL+qd/+idoF8jHQ8+gU0oppZRS3xsRoWfPnvHJyUlmrR157+fMvPDen8UYr8bj8eP5fP748ePHN2dnZ1enp6enRVHk1lpDRLr66gDtn13ZNA3W6zVub29xd3eHzWaDtm13JegP110NByQO+SDErvODqAs/RGCl6/uwMXaTHM6B6qab/KgqpKpC3JZIVbf2KtY1YtMA3oGcA4XQrb0KAeM+/MhTAkPAH/LGHoHIjMAGnhmJGcTcldkTdz9ja8E2A1kLNhZkDNhwV/kBIEEQRZCINPRQSqk/guGxxH4XyGB4jDGsxhqNRphMJphOpyAihBDQNA2cc4gx7v6MPlw9DP3PkpiZrbVMRCnG6MuybMuydN57z8w+hBCzLHMAvPc+/dVf/VX8t3/7Nzx79oy++OKLw32Q+gnRAEQppZRSSn1f6NmzZwzAfP3114VzbsLMJyGEZUrpPMZ4PR6Pb+bz+aPr6+vrs7Ozs9lsNrfWWg0/DldKCSEEVFWFzWaDu7s73N/fY7Vaoa7rXfgB4FsByEEbDsgAIJHd5IcFgVOCCRE2BBjnYFoHqusu7Nhuu0tVIVVd+CFNjdS2gPegEMAhwISALEaMYkQuCVaSdn58DyIxAlEXgBCBQbAisAAMETjLQcb2QUgXgkjf9ZGkm/6I6MIQGf5L1P8alVLqD/a+Eyn2X99fi2WtRZ7nsNbuHrus1+tdALI/IaIOAvUrsdgYwyISm6YJ9/f3brPZ+KZpAoBARD6l5AC4lFIoiiJ+/vnnuLy8xA9/+ENoCPLh6QospZRSSin1vXjx4gV9+eWX5kc/+lFmjClEZOy9nwM4iTEuReTce3/Wtu2pc24cY9THqkcgxoi6rvHmzRvc3t7i/v4eVV3Be/+taY/3XT9YD85AZWYYEVBKMCmBUwR5DzgHNF2xuVQVYlXBVxWkn/xITQ3pVytxCECMoOEiqVt5deDfyo+LAJKAmLq+jxiR1RWytoUNASkvgCwD8hycZRBjYKkLCmNmETmDBSERdsHI0AOiP0allPrD7E96DK/vv29YeeW9x/39PZxzu5DDe4+TkxOcn5/jyZMnu6BEHZ4Yo3XOjeu6Pm3btmzbtkkpNVmWtSJSpZSa+XweYowxhOA+++yz8NOf/hQiIroO68PSf5FKKaWUUur7QAD48ePHdrvd5lmWjZxzExGZMfNJURSnxpjldDpdjsfjhTFmTESme76gZzcfmmHtVQgBdV1js9lgtV7hfnWP9WaN4MNulcT+nwGwmwY59NVXwLf7P9BPglBKoBgB74HWIbVNN+XRNIhNg9S2/UuH1DrAeVCIkBC6CZCUYFOCTQIS7f34PpEIOHUrzEgEJgZk/VozZkaaz4HxBDKqgSwDWwsQgfoVZYYZ1hpE4t0USOi7QGgIBvX/TKWU+r297/HmsM5qeF9KabfySkQQQoBzDs45WGtxcXHxTl+ZOij9MIgp8jyfF0VxGmNsiKgKIdQish2Px1Xbtm48Hof1eg0AuLq6kpcvX3ZbLPVchQ9GAxCllFJKKfV94bZtrTGmCCFMRGQmInNr7WI0Gi1ms9lyuVyeLhaLk9FoNDLGWA0/DtPQ+TGEH+v1GqvVCpvNBlVVAQCoP/z/sJz0fdcPzv5ZqP0FScDSHUBHSkAYSrQd0LRITYvYtkhti9C2SM4jOgdx3dorihEcIzglZEMAIt1Bdf1X9v0h6XtcUoSk2K2/SgmGCMgyUNNA6hqoa4i1IGu74l0msGGwMV0IwrIrRmcixOGAm/6fqZRS/2dDEfp+/8fQRea93z2OGcKPLMuwWCwQQtAA5IAZY0ye58V0Op177xtmbuq6LmOMVUppE2PcGmNaZvbW2nR7eysA4t3dnYhI0uc1H44GIEoppZRS6k+NXrx4QScnJ8Y5lxdFMQYwJaI5gJOiKBanp6fLm5ub5eXl5WKxWMy67vNC++oO1DD5cXd3h9vbW6zXa2y3W4QQugP/e9kGEb3TAXJM3l3H0R08p34NFmKEBN9PeDgk5xCdQ/Qe0QdE75FCAFLs1maJgFJ3sL2QhJF0L61oAPJ9YnQ/gzG6X3MWgZEEpG5CJ7UtUlMDVQU2BmIMhAlggjEMm2WIKcHCdH0g/c+PiZBE9NRSpZT6IximTIf74YeByMOQw1oLY4wWoB8wIqIsy8x8Pi8A0HQ6be/v75vXr19vt9ttGUJYE1EJwImIjzGGxWIRV6tV+PzzzwXd+Sx6N/2BaACilFJKKaX+lOjFixcEgBeLhXXOFc65aYzxREROQwhLY8xyPB6fXl5eLh49ejQ/OTmZ5nnOxhijTyIPx7D2KsaIqq6w2W5we3uLN7dvsNlsEML7117t934cExEB92EQEYEE3WTIMAESE/4fe3eSHMmV3A387/7ei4gcASSAmr4m25rWkslI7VpLyVoLXaF0DZnpAiqeQUeQmRaiTqBV9QF6J/ZCppUGssWakMgp4g3u3yIis7KKbInsrmIBVf4zS8NQIJhAIDMj3v+5O3IZgpAMSekQfkjO0FIgpbwMS4r0LZdUUQ0hSLVvqfWuf9gPCAHwUPC+ldtQgaOi/fFqW2CzAfkAAQAmwDHADPIeXAV47yDq4QEUBbLo4fvY6ooxxrw5xwPQj8MQoA899ucp+wqRGCPatkVVVYdh6DYQ/f1ARHDOufF4TFVVuaqqZt77mFLaEVG32+22IYQOQO66LldVlVarVfHe51KKPH78uKBvg2XeAQtAjDHGGGPM20IPHz7kr776iv/0T/+UVTWklBpVnajqvJRyqqqnRHTivZ+PRqPpdDodDzurzHtm3y5iu+3Dj+VyieX1EtfX19hut6/umqR+QRh4GYIcV0N8cLRvd/St4ayqUBluRSBF+iqAoU0HVAEZhpwP4QmjD0G8Av4DC5VuAtpXbLwWU6hqP6OlbUF+DXIOCkC8A5wDggfVAZxquNDPbxFVOAIcEfajPwgfXlhojDE/huNzEGZ+pUoE6Ktb1+s1qqoCM2M8HiOEYAHI+4Occ+Sc46qqPBGNRGS23W47Zo51Xe+IqHXOxZxzp6o7733sui6enZ3lr776iofZhvYi/Q5YAGKMMcYYY94GevToEd2/f583m42fTCZ+u902XddNcs4nMcbTGONZjPGs67qTnPMk51ypql0lvqdSStjudnj69Cmuln3wsdn0ba/2ky5UFQSCQl9ZxP1Qg49D6EPD7wd9EAIaKgKcAzkHeA+EAOdDHyQNbThAQ/UIhsXxD/PXeDtIAaUEt1mDVVFEhgCkP7ZaVUBVgesI9gE+BCg7FAKSKnjfOW4IWGx1xRhj3qzjjRj7ig9mhnMOIoL1eo2vv/4au90OXdfh4uIC8/kc3tvS6/vIORem0+n47t2757PZTDebTV6v13m32+WUUowxbr33nXOu++abbzKADCAPf0f2Mv0js0ehMcYYY4x54/Ztr6qqcr5XqeoIwCTnPAdw6r0/I6KzEMIJM88A1AAsAHmP7NteiQi6rsNqtcLzFy/w4sWLw8yPUspRRQMg+u3uAB/ajnZFP9OBjj5WAvpGR+irQZhBAloCiQAAIABJREFUrh+SDedAzoOd62/MUO6Hth4nH3R0MzcLqYJzAu0URQUqBcU5aKigVQBVNWg0AmKCqzOQC4QLvHPwRJAhADk8emweiDHGvBGvn4McV2MeByDb7Q5t2yHGCACo6xre+8PX7KtGzPvBe++IaOS9903T6L4dVtd1u67rtsy8BLAtpezquo7OOf/rX/86/+IXv9j3e7WX6R+RDZY0xhhjjDFvGv3lX/6lWywWLoRQ5ZxrERm1bTvf7XbnpZS7zrm7VVXdPTk5uXt+fn6xWCxOLy4uJicnJ3Vd17ZJ5z2x74e92+1wfX2Nqxcv8PTpU6xWK2y328MQ0eMFgdd7bH9o4ccBUb+b/1DBQWD0CSFJAYuAi4BzBhcBlYwSIyQmaM5AztCcwVLApYBV4UVRqaBRRQDg7Nr7RukH3Jf+rSpUCcoMZQYHDwoBVNegEPqqH+cgTCjUh2KCISzDh1s1ZYwxb9rx8+l3vb8fip5zRte1h3lmx6HHfhaItcN6fxARMbMPIQQiopSSrNfrvN1u4263iwB2qtoRUZdSKk3T5FJK+Zd/+Rf82Z/9mT5+/NhOwn5EdnFpjDHGGGPeqEePHtGnn37Kbdt6Va1EpOm6blxKmYrILKU0b5rm5OTk5PTBgwen5+fn87Ozs9nZ2VkVQrANOu+RnDM2mw2urq5wdXWF5fU1drvdoerjlbkfR3M+ROSV3tof2mIuDeEH6GXFhw47+gUAgeD4aDZECCAf4EIF9h7sPNT1C+RK3FeFiAwzIqh/a5fdN8txy7dSQDHCbTcg34cc2jTAeAK0HWiUwKmAfYEjgiMHR/3fxr4CZB+EHIaDGGOM+b191znJfvj58awy5/yhHdZvf/s/6LoO2+0Od+5cWjus9w8NfwsEwKlqPbT0nccYT6qqmhHRFMDKe9/Vdd0CiB999JGenZ3ZMPQfmT3yjDHGGGPMG/Xpp5/SZrPhGKOPMdbM3BDRWESmAOaqOvfez6fT6fzevXsnd+7cmZ2cnIybpnEhBNsad8vtFwFEBG3bYrVa4enTp1gul1iv10g5HwKO/U7I16s9PuTw45gehyDo55kzAGXqb44BH0BV6EOQEMAhgL2HOgfdzwnJ+6CJXva/skERNxapgnKGa3f9rBfvUWZb6K4FxQTtIrhOcCGAmeAcwylQQHBDeFYwHOIP+PFjjDFv0nF16t7+PKU/p3EACKX07bBiTOi6DjEm1HWNEAJCCIfznw/5/OZ9IyJORCoAEyKaMfOJqs4BLEVkGkJoRWSXUoqlFLm8vCz/1/c0b5YFIMYYY4wx5o36zW9+Q5988ombzWbh6uqqyTlPRGQO4CTnfFJKmQOYOedm0+l0PJvNRrPZrB4uBu1q8JYrpQxtIDpcX19juVxiuVxitVqhbVsAAB21gVBVqMgriwrHQcgH66gFlmo//FwJKBiGrx7CjwJNAVRX4LoGVxXI97NB2AeAI8AO4AJiAsp+CoilHzdVH/4JJGdIStCug3YRGjto24K6BhQjOAR47+BE4Zn7OSDHgRmGI/2htpEzxpg37PXzkv3HzjkQ9ZWWpQhKKei6eAhIptPpoVqkaZrDfBDzfiAi9t5XTdNMxuPxXETWOecTEblm5hUR7Zh5t1gsOhHJ//Ef/5Hf9X3+0NijzRhjjDHGvEkEgJ89exacc42qjolorqqLUsq5iJznnE9zznMRGRNRzczee2+VH++JlBJWqxWWy+Wh9dVms0FK6WVFx77iYwg+9jfAFmtfcbTbVFSHWSD9wrayg3iBVgFcGmjOoLZ9GYJUFUrXQX3o/60wQPuh6LD84wZTAIUIkRiFCGWoCOEugtsW1LZAXQO+H3wfHAPMUMdQ9EGZiMKiLmOM+XEcb9xwjg/tsXLOWK/X+Oqrr7DbbbFer3F5eYGzszMLQN4j3ntumqY+Pz+fNk0Tp9Npu16vF7vdbt113aaUElNKbdd1saqqdHl5Gd/1ff7Q2KPNGGOMMca8MaqKv/3bv3XT6dSnlOqqqiYxxn0AsiCiM+fcydATt1FVb1Uf74fjtlfX19f45ptvcHV1he12i5zzK3M/dPj6w1sLP34nOe43PtyECMIEcQ7FB3ClQF2BhvDD1TWk6wDvId5BHYOY+wqQfSssc2MpqA9AnENkhpCDF4GLEb5tQW0H1C2oquCqgCChf/wpIAQIhr8PsQ4bxhjzNh23wDq2H4Cuqui6Dt988w222y222x2cc2iaBlVdg1+fh2ZuJWZ24/E4DEFIapqmFZHTnPP1drtde+93pZRNSmm32Wx2RNSqKhHZRLYfiw2ZNMYYY4wxbwoRkfvoo4+qruvGIYRZjHGRUjpX1QsAd6qqujMejy8uLi5Oz8/P53fv3h1Pp9Oqrms7L73Fcs6IMWK32+Hq6govXrzAs2fPsF6vD22vgJetIvaX+a9Xf5hve+V3pi939TMzeHifAFARaMrQGIGcDzcqApQCKgVOBPVwC6pw9nu/kYQJhRmdc4ghoIQKCGFoeVYBzIB3/ZwXx8O8F+qHoOswDH0fMAI2BN0YY96Cw+vza7NBXs4E6QOQUgratkWMCSKCEAL8UMGnImBmOGenwbfZcLzZe++ISEQkr9fr3WaziZvNJqpqIqLOe9+1bRtjjPG3v/1t/tnPfobHjx+/67v/QbAKEGOMMcYY8ybQP/3TP/Fvf/tbR0SBmeuu68allGnOeQ7gdDQanc7n89OTk5OTxWIxPz8/H08mk2Dtr243VUVKCev1GsvlEi9evMByuTy0vdoPPD/++tff/9CHnX8fiqPh8Ez9QrdjFHFgJ4D30KpfIOeq6lsk1TU0RpAP0JDBpYBy7n/X9uu+0Q7VUaIoJYNzhqSIstsBVQXdVaAQIK4PQgCAKgEPi2qOqZ8Jgpd/O2KBlzHGvFG/aybI8Mx7+FhEEFPEarXGk6dPQUToYsRiscDJfA7vvZ0H3WI0AADnXGDmOuc8TSnNU0onIrJh5uu2bdfMvK7rugLg79+/X1S1DN/DXqTfIgtAjDHGGGPMH4oePnzIANzp6an/7W9/W+ecR6WUSUppWkqZq+rpfD4/PT09Pfv4449PLy8vZycnJ+PpdOpDCBaA3GIighgjlsslvv7660Pbq/3Mj+Ndja+3uxIRAB/4sPMfQPFyyLVAUYjBHigiUO9AIQBVANc1KEbQEIBoTpCSwTmBHFsbrJuuTz/6m/QVPJISStcB7Q4SAtg5ELs+2HDcV3xIH3qRCsg5kHNgftly7vVdysYYY96M76oC2b91ziGE0FeCdC3+53/+B7vdFqv1CgDQNA3Gk4m9Kr8nVJVLKaGUMk4pzWKMp1VVbbquWxLR2jl33XXdZjKZ7P74j/8Yv/71r/GLX/yiDK/T9iL9llgAYowxxhhj/hD08OFD/uyzz9yTJ08qVa1LKeMY41REZiGE0+l0elbX9fnFxcX5/fv3T+/evTs7OzsbTSaTyntPzGzXfLeYqiLnjK7rsF6vsV6v0XUdnHMvZ1e8NuPjOPiwBdkfpg8/ACaCMJBEAceA96AQwM0IGhM4Z1CMQIzQoQ1ZEEUQgVMF2WjsG4sAOFV4FXgpQErQ2KG0HuIDmPve8v3jS0FMEBGoCKAA1RWYCN45ZPShmQAgVcAec8YY81bsz2lentu8bIXlnOvPl0rBbrc7bBDZ7XbIKfWBt20GeS8QETvnqtFoNJ3NZqciEkVkW0pZdV23CSFcj8fjjYjsRqMRnZ+fx30IAtjJ2dtiAYgxxhhjjPl90aNHj+irr75iAL7rusp7PxKRMYBpjHE+n89PTk9Pz87Ozs4Xi8Xi8vLy5PT0tJlMJsHmfrwfjts75JyRcz5Ueuwv/Et5OYzZFl9/f3r0VoB+wYQZWRTqGL4K0KoCNQ0oJdBoBOy2cN6BVRGkoMoZTqVfDDc3EkHBCgQRaCkgzsgpQWKEdB3EO4AZPDy+yDlI3+cKGCo/yDmwV/A+6tq3T3vHP5sxxrzPjkOQfQBCRPDeH1oS5pxRSkHOBUXE2hO+Z5iZQwjVfD6fEFEMIcTNZrPebrfLruuWzDxLKa3Ozs42zKz//d//rXfv3tXHjx+r9pPR7Q/iLbAAxBhjjDHG/CG4rmsG4ImoTimNSymzruvmqjpvmub08vJy8dFHH12cnp4u5vP5bDweV86mPb5X9i0evPcIIbzS+up4N+Tr4YeFIT/QfofosKMfDJAC5B1IPIr3/e7/XPcBSEpwVQVPhJATfOwQUoSTArbf/Y1FABwUtQi4ZDARdimhcIt0qPwYdhbj8CcBDAPR4R1c8IAqHPp/VBHwUfWH2m5jY4x5K47ngPTPz3SoAFHVw7lSCAGOHawN6PvFOcej0SgsFovpaDSS0WhUnjx5ss45v9jtdnMRmTHzNOe8YWZlZlkul+XJkyf6+eefC6wK5K2wAMQYY4wxxvxeHj16RAD4448/9pvNplqv12NVnQ1Dz09KKafe+5PRaDSfz+ez09PT8Xg8brz3bG2vbrf9/I6cM2KM2G636LruMPCcuR/rQjS05jkKP/ZfY+HH72GY/6HAt3eMEoGcg4YArWpQ3QcgVNegqoKrAtwwILsPP6QPVMyNQ0AfbKCfAyJS4EoGsoOkBO3a/ngT9V/LDBoqQaiqgFSBcoHbhx0YFuRUQbCVFWOMeZteVoBgqADZF+g5KBSqAc4xVBVd12GzXmPVNKjrGt77V1qImttnqAABMxMzj0RkslqtJvtrpBDCHMBqGIxevPf5xYsX5fLyUj799NP9kDZ7qX7DLAAxxhhjjDG/j/0aHZdSvPe+JqJJSulEVc9yzgsRWZRSToloXtf1uK7rpq7r8K7vuPnD7ed+bLdbrFYrXF9fY7PZHFpd/a7ZHzaI+c2Qo4VsBUEIIMeQ4KGlghYBSgZyBo3GoPEEmEyBlIBSoO0OlDOGRlrmphmObz8LROCFQKVAU4ZQBwEd9UPTvhWWY3DwcE3Tt0Ar+SjwIBRVlNcG9Nqj0Bhj3rzj8KI/7wEAAjPBwR2+ppSM6+USVfBQVZycnGA6nR4qRsztRD3HzE5EqrZtGwATALNSygkRnTLzZpgLkne7XfLe5xhjvry8zO/6/r+vLAAxxhhjjDE/2L76YzKZuM1mE5xzTc55KiInKaV9+HGWc57HGMellKCq/K7vt3kzVBUxRlxfX+Pp06eHAGRfBfJdba9ef2v+QMPvVw4fEoT7EISyB1cVtK6g4zHKbIYUIxQEFUWlAlUBlf/1/2BuAkVfqVMKQBmaGEqxP+5DiEGO4YKHqytwjOCU4ESAIiBRCA9pNYbFONjWUmOM+TEcb/ogor4VIb+s/nj67Cl27Q673Q6llEN7LPN+UFVSVVdKqXPOY1WdicjJUP2xYeY2hLBLKbWlFDebzei4gsi8ORaAGGOMMcaYH+TRo0f8y1/+kn/1q1/5nHMFoCmljGKMM1U99d6f1XW9cM4tZrPZyXg8HjvnAvr1N3NLHbe96roOq9UKy+USV1dXWK1WiDGilPJKi6vvupk34+VCtkIJUCLoMAybqwDJGVzXkKYBTaeQnFFKhosdZLcFUfeufwTzvfRtsKAKKgKiAuQMJYIQQamfAYOqAncR6LqX81+Gx6MIwQH91+Nl+zSCzQIxxpgfw6stsfpzpFIKttstcu43/VdVdZijNhqN+hkh1g7rViMids75qqqayWQyyznvqqraMvMuxrghoi2Ajfd+d3p6Glerlfviiy8EgG1RecPsItQYY4wxxnxvqkoA+Fe/+pVfLBa+67oaQJNSmuacZ6WUE+/92Xw+P7t///7ZxcXFyWw2m1RVFXg/GMLcSiKClBI2mw2WyyVevHiB5XKJ6+tr7HY7xBhfmfexD0ws/Hh7FDhMwFYiKBPEMYpzkBAgVQVtamjTQKfT/tY0QBUAZw/HW0MBEgWJDK2wEjQlSIzQGCFdN9zaPgCJEZwyXC7glOFFwTrciOCG2SH7hThjjDFvx+vzQJi5n9sEQEpBivFwXvX8+XM8efIEz549w/X1NVJKELFWlbcZEbH33o/H4/HJyclssVicjsfjMyI6SymdlFKmIjIWkXq73YYYo/vkk094uN4yb5BVgBhjjDHGmO+L/vqv/5r/4i/+wu12u9B1XVPX9Xi73c5KKfMY46lz7qxpmrN79+6df/TRR5eXl5dnp6en08lkUoUQbMX1FhMR7HY7PHv27HBxvt1uD8HH6z2v9xftxwGILba+HTL8bgWAOAZ7Bw0OWgLQNEDOQCngZtQPRXce/f5/c1uQKkgVLAImgpTcF25kNwQhHdD1N+o6cNfBxQhyDPWMwAxlhiggIDimvhLEZvIYY8xbcxx+7J9r922wjsUY8T/ffIP1ZoOr5RL37t6Fc+5wM7eTc45Ho1F1cXExHY/Hutls+Pr6Oq9Wq7jdbtequmLmVVVV21JKIqL09ddf6+PHj1VVCxHZC/QbYgGIMcYYY4z53j777DPqus6XUqqU0khEJgDmo9HoZDQanXnvzy8uLs7v3r17eu/evflisZiMx+M6hOCsAuT22bdoOG57dXV1hefPn2O1WqGU8q3qDgs/fjz79kV0aG2EQwhSnAN7DwmhH4ydC3Q0gjYjSN2A6gaSIqgU0NBiydxMhL56ww8D0YUAKX1LK0kJ5N2h7RW6rp8DMoQgcNwvoAUPN1R/gAgFCiXqW2tZCGKMMW/V68+x+0HnRDS0KhRsNhu0bYsUI7z3mEwmYGZrh3WL7StAJpMJee+lqipV1VZEWhFZiciylHKVc14751pV7ZqmKQDkiy++UPSndfYC/QZYAGKMMcYYY76X/eDzUopX1UpVGxGZeO/no9HobDwen08mk4vLy8vz8/Pzs8ViMZ3P500IoXrX9938fkopSClht9thvV7j+fPnWC6XWK1W2O12AHC4IN9f3Fv48SN6reoGTBAFihDIO4h4aBWgRaCjAhqPoZMJZDoFuhaaE7hrwTn3IYi5cQgAQ+GhCCooIIigD0GEoCVDUwJSAmIExwi0Laht+wDEe7APYO6H7zrnABrGiqAPUSz8MsaYH9fre4IkZ8SuQxGBlIKqqjAejaCqODk5wXQ6RV3XVg1yyzAzAXADOOcQY4wiEolo3XXdi67rnqvqtYjs6rpunXO5lFI++eSToqpi59Bvhj1yjDHGGGPM93J5ecl37tzxzNyklMZENC+lnFVVdX5+fn7vo48++ulPf/rTj+/fv3/3/Pz8bDqdjrz3NvvjFtuHH0+fPsU333yDZ8+eYb1eI8b4SrBxvLPx+HN20fYj2A+xHkIoQr9oToph7gPgqL/wo9LPkJCjyh0WOcyWMDfQvn0KXg7wVOqno8pw3EEEdg4+BPgQ4KoKzvs+nHQOcA7qHMAMMB+2kioNFVsWgBhjzI9mP39pPxPk+Lxpfz5VSkGM8XC+1TQNqqqyAOR2UyIi5xyHELiu6+Kc24rIJue8U9VERLmu61xKKcvlsvzjP/6jPH782F6k3wCrADHGGGOMMd/LZ599Ruv12k2n0wCg6bpuAmAuIvsQ5OLevXuX8/l8MRqNJt774JyzFfBbTFURY8T19TWePXuGq6ur31nV8XobLADfmg1i3oJ99c2wEC7D54gZzntIpX1bLAV4miExAl0HEYGDwpXSByAigIi1w7phCEN4Be0DEJW+ykcBlQIqhFIKOGdwjP0A9LYFtltoCGDvwd7DOe4DE2YIM5T6aiElAqlafw1jjHnL9udGr58X7dthee8PrUfX6zW6rkMc2mGdnZ1hMpm8i7tt3pChHVYYrpEQQtiKyGKz2ZzlnJellNZ733ZdF6uqSnVdd59++qmdRL8hFoAYY4wxxpjv5auvvqIHDx44733ouq4monHOeaaqJ865k6ZpTmez2Xw6nU5DCM27vr/mD7ef/9G2LdbrNdbrNYaLtu+s/gBetsACvn2Rb96SYQYI0FcG0DBgVQBoGAIQACU30MkYaGegFIEUUXY7UMlAyeBhWLq1w7pBhqoeB4AJUCiKAkX281/66h0qBYgR2raQ3Q6oKqCqoCGAqgouBKj30JThgocM80AEw0BefPuxbIwx5s35XedE+6qOfQAiIogxous6hBCw2+2Qc7bn6FuOiJiImJm9c05VdRZCmAGYA5iXUjYppU0IoY0xtiEEf3l5md71/X5fWABijDHGGGO+D6rrmtu2dd77qpTSqOokpTTLOc+7rpullJpSike/adm8B45bMzDzKx8fz/04bttgA5XfHVU9LGYLAYUIhR3Y99UDlANQV6CmAY1GwHSK0nUA+kVwv92Cu7avBjE3kgNQDY8vJwKmglYctBQg55chSFWheA/yHhRCPwvEcT8HBIB4B2HGcX9Ce+waY8yPa/+8u2+J5ZxDCOFwXhVCgPfeNpS8Z1SVVNXnnEciMhWRuYhsVHUTY2y997uU0vrf/u3f7MC/IRaAGGOMMcaY/ws9fPiQz8/PXdd1vpRSq+qImSej0Wg+Go1OQghzIhoRUd+txdxa+4tuEUFKCTlnAC8DkP1Il+9qeXX81i7W34HDTn5AQX0IwgRGP6geVYCvK7imBsZjICWUmKCq/WJ6yX1liLmR9nNAKiicAqz9NHSRgpwSKCVo10HbDtltAefhfACFClRVIO/hmFFU+/kwwfWt0oa5IAq8bKlmjDHmrTg+RzpuFXo8Mm//PHzcFiulhJTStzakmFuJRMSXUpqc8yyldFJK2arqWlW3McZ1KSVUVeUAZMA6Vf6hbHqOMcYYY4z539CjR4+cc86Px+NGVScicuq9Px+Px3fPzs4eLBaLB5eXl3cvLy/P5vP5tK7ryjlng89vKRE5tL1arVZYrVZYLpfYbrevXHgDr1Z+WPhxQ6gO40Do5XEYJqOTAlwKWEo/EF21/wcRkBRwjHBd17fCMjcP0SEEYfTHE6B+jgcTmB2IGMT9DfvZMM6Bvet7aO3ngAxt0nT/9vX/1/6/NcYY80YdtxD9rnkgx5W2VVWhaRrUdQ3n3GFw+vG5mLl9RERijHG1WrXL5TJut9tcSsnMHIkoElGbc96enp7Gf/iHfyhERI8fP37Xd/tWswDEGGOMMcb8Tg8fPnR/8id/4sfjcUVEE+fctG3bxWg0ulgsFvc//vjjn/zkJz/5yb179+4sFouT6XTahBA821XZrbUPP168eIHnz5/j2bNnWK1WiDG+slNx37bh9aGeFn68Y68vpuDouIiAVMBFwKog1X4AeukHaLvdDq5twclaTt90h8fbcGOi4Z0h1EC/XZSY++DDOSheHYIOZqhjKPfvH33zl1Ug9ng2xpi34vX2V69//nizyb4id98WK4RwmB1ibh8RkbZt8/X1dXzx4kXa7XYp55yccx0zd0S0q+t6MxqNUoyx/PSnP6W/+qu/whdffPGu7/qtZY8WY4wxxhjzu/Df/M3fuO12G5i5UdVpSmleSjkfjUYXd+7cefDRRx/95MGDB/9vsVhczGazSQghOOeYbBX81hERlFIOA8+fPn2KZ8+e4erqCm3bHlphvc7a5dw8xw++Vx6JqnDDjUUPIQjnAooRbrsDty0oZQxlJC+/yXCjo/fNOzRUgxAUDsPhIEIhghC/bGdFAJwDOdeHHM71t+F9dQwdPt6HJophAe6d/XDGGPNh+K4KkP3b/SaTlBJ2ux1KKSAi1HX9rQDETrtvl1KKxhjLarXKm80m73a7AiARUcfMrXNu65xbV1XV3bt3r4QQ0DQNHjx4oFYJ8vuxAMQYY4wxxnwXevjwIY9GI++cq7z345TSXEROYozndV3fWSwW9x48ePD/Li4u7s3n85MQQnMUftiV2C2y7y292+0OLa+eP3+O5XKJzWYDORqK/V2Dko93MZob4CigoOFj2rdPEgUr+vADfQUIUgZiAnctNHaQklGYkYlRqG+XVPCyquDwfc2781o7LBBBiJCG4yXAUB5CfRXIa8EHnAN8f1PnAGL0cYr2x9haYBljzI/iuNrju+ScEWM/n4uIDkPR9/+NtcO6fVRVY4zadZ3EGBWAOOcSM7ci0hLRZjKZrOq67qqqytfX1zqbzXSxWOBnP/sZHj9+bHsUfiAbgm6MMcYYY74LnZ2dMQDftm2dUhqXUqY557mInIjITESmRNQwc8XM3uZ+3F45Z+x2u0PocXV1hfV6ja7rXvm64/DjuP3V/t/MzaJEkP3xAgAiOO8hlUCkAatCcgaNO+h0Cp3NQV2EgqApQXMGSgFKBonAiSCoIKjCUs537JXH3hBoFQHlDHCEAhAolBkIAfAe6hyc90BVgUIA1xW8CFQU5AmqAkH/t1LQH19bYTHGmLfr+Nzqu1ph7T/XdR2urq6gqthut9jtdri4uAARWTusW4aIqK5rP5/PR8wsk8kkbzab3Wq1WnZdN8s5T2OMk9lstlqv11FEsN1ucefOHf3000+HAW72Ev1DWABijDHGGGNeRw8fPqT//M//5PF47Kuqqsbj8SjnPB2qQGY551lKaZJSqlW13zpsbh1VhYggxoj1eo0nT57g6uoK19fXh5ZYx8M6v+sGWPhxE+138e9DEAKgzCgskKqCaN/2jGIEjRpgPEaezqBdhKhCY4R0HbTr+sHaOSGAoAI4LdZK4KZRBaQAeV/901fsFOdAVdXfug7atkDTgOq6D0tyga+0b48G9MPR0YdnZZj5Y23ujDHmx3H8fPt6i6tSCtbrNdq2PbTEGo/HaJrmXdxV8wdgZgohuPl8Xtd1jaZpsvd+07bttOu6iapOVHXcdd1IVeNut9O6rvX58+fl8vJSrOr6h7MAxBhjjDHGfMtnn31GX375JTvnPDNX2+12XEqZq+pJSukkxjiLMU5yzlUpxdZCb6GcM1JK6LoOq9UKV1dXh/Bju93COQdmfiUA2b+1yo9bYj/HYThGAkDYIUNBzgOhAoUKVDdAM4KOR9B2gpILhHcoqlARQAGnCmiCB0GGVkl25G8GAkDDbJcgAskZIEamvpJHug7cttC6hlYVXIxA7ED2nICGAAAgAElEQVQxgusKVCpABAWKcpgt0rfW2j/SLQIxxpi37/XQ+XgQeinlULFLRJjNZui6DqWUd3V3ze9pqNphZibnnAKot9vtiIgmIjItpcyGavuVqqYQggCQxWKRU0rl888/twqQH8jaFBhjjDHGmFc8evSIvvzyS768vHSllJBSalJK05TSSdd1Zznnk5TSPMY4zjnXqupU1dZCb5mcMzabDZ4+fYonT57gyZMn2Gw26LoOIgIReSX0eP2t7T67HVT1MLujD0AImRnZO+QQkENAqSqUukZuRsijEcpohFRVyKFCch7ZOSTazwQhqB33G4egcCqopKCWglAyXM5wpYBSgsYIdBHaRaDr4GKCixEuJbiU4HOGE+1nxKBfKNjPjbHHuTHG/HhomNu1f985d9iUAuBQobsPPqxK71aiIfxg771j5gCgFpFRznlSSpnlnE9jjCellKmqjtq2rXa7nfvmm2/47/7u7971/b91rALEGGOMMca8jieTCc9mM7derysRGZVSZqWUUxFZ5JxPq6qap5QOFSAWgNw+OWesVit8/fXXh5kfOWeo6mHAJvDt1leALYjeKsdzW0D9bAcG4BjqXT8LIgSgCqC6htYNpO5QYoT4CHEOxNy30mKGih37m4gBBFU4CFgIJAUijFIKpBRQytAYQTH2bbDqGtTUoK4GVzXIZ3jnUJxD1v4xzkP7NN23UHvXP6QxxnxAjs/D9kPP92GI9x7OuVeGoZvbS0S4lBJyzk0pZaKqcxE5K6Vscs7RORdLKSmE0J2eniZY6+EfzAIQY4wxxhgDABhCDPr7v/97B8Cv1+vae9+IyDilNPfen1RVdVrX9dnZ2dnJxcXFdDQaNd57Zwvit08pBV3XYbPZYLVaYbPZwHsPZn6l5QLQ7zY8/tjcMkMIohjmgKgOk7MJ5Bw4BHBdA00DNDWkrYEUISlCYgKVApSCooLEjKgMFsBDDq2SYH8b79R+EBOrQlWAIhAqKLlvgUXMYO8Ax3DNEH7s+vBDqwrsGBwCHBECOxAIBXRYYinazwmBPdcbY8xb9/pg9OMQxHsPgBBjwmq1RlVVAIC6rg/BiLlVyDnn6rquZ7PZlIhOcs4b7/1aVbcppS7n3KaUEhG1zBy/+OKLgr6w106+vicLQIwxxhhjDADg888/p/v377u6rl1d1+H6+rp2zjWllLGqTpxzs/F4PL979+7JnTt35vfv35+enp7WVVU5sgTk1tkPQE8pIaWEnPMh/NhfbB9XfRyHH9b+6hYa5oH04QdA3Le0csFDvYeGCjxUgOgoQmIE6r5lkuYMGtptJBZEURD1V91e5TAzwrwj+0Wy4eZFoSiQApTYV3GQ9OskxASMR0BTA3UzVINUfRC232HMDGWFDsdYMSzAvbuf0BhjPhjftdlk3xZrf56mKmjbFs+fPwPQzwc5PT3FeDy2AOSWISIKIbjxeFwvFotZ0zTdbrfbxRg3qrre7XZb59xGRNqU0ialFABkVc3Dubi9PH8P9qgwxhhjjDFQVfrVr37lzs/P/dOnTysRqUMI467rTnLOi5zzvdFodG+xWNz55JNPzj/55JPFT37yk/nZ2Vk1Ho+9954tBLld2rbFer3GcrlE13XIOSOE8Mrgc+DVuR/HuxDN7dQfOgIp+oVzEUAEpAKUAuQCyRlaCkpKQCkgEWgRQBWEl9UkBMCrHqoPzA1BAGl/se9VUJWCkNNwrKgfhu4DEALgHMg7wDmo84DzUMcgZggAMB9CEGOMMW/fd51jHX9ufy5WSsZu16LrInLOaJoGdV0fKkLMrULe+/0mNDjnJKWUuq7rYoxRVVsAXSklxhiT976s12t58OCBPn78+F3f91vBKkCMMcYYYww+//xzAsDb7daPx+MqxtiklMbT6XQymUxmInJ6dnZ2enFxcfrgwYPZnTt3xufn53UIwXnvyfoP3z6v7ybcH8PXZ38cs/DjdtsPQqf9kjb3bbCwnwVS18CoAeUMpAiOI0iMQwusDKigqCKrhwdQoBAVa391w/SBlIJF+sew9OFWIUJhhq7GoBAgIYC8B6oKCFXfCs37vr0KCbxjqPbfT2wKiDHGvDPH7bD2AUiMCTGmvu0hFJPJBEQEEUFVVQghWDXILTAMuue6rr1zrvHeTwG0OecdM6+7rtvEGJequs45r4iorqoqrVar9Mtf/lJVtdi5+f/NHgnGGGOMMQaXl5f885//PIQQ6mHo+STnPJ9MJuenp6d37969+9MHDx589ODBg3sPHjyYn5+fj6fTae29Z2a2Dji3UIwR6/Ua19fXaNsWOefDQM3jFljm/ULf9Vb7ioH+/X7Wg5YCLaWvDjlUiejhxlA4EVSqcAqwLY7fKP2TsoJVwSpgEdB+pMfQv4wAwDHEecAPN+f7ihBmKAggggAQKNTaYBljzI9ify723R/TUMDZtzEtpUCkAOg/V0o5zArp54WYG46IiJiZnXPsnDv+uBBRVtVtzrnrum4nIomZcwghP3nyRP75n/9ZHz9+bC/P/wd7JBhjjDHGGHz22Wd0cXHBOWf/9OnTupQyEpHJZDKZX15ent2/f/9isVhczmazxWQyaeq6Drbb6Pb7rgqQ12d/7D9n3g/71lUyHFIiAjuHEjwINXhoeUUxgmIEUgJyAZeXQYiUApUCZQbKu/xpzA9BpYC7Dv56CRJBEUF2DqgbyGgEqmu4ugZKgTqGHwIPByADfQu0o8G8xhhj3q7Xn3P7aoGXlbrOOYgUbLdbfP3111iv11itVgCAqqrQNM07ud/m90bOuTAej6feezcajbqmabZE9CSldKWqE+/9pqqq1nsfLi8v86effmoXZN+DBSDGGGOMMQb379+nr776yldVVYlIo6pjANP94PPz8/P5YrGYTafTiffeOaupv5X2OwNLKdjtdkgpQUQAAMdtzGyR8/3WD7Ueij2YIU7B6vth2XXVz/0Yj8ApQlPqW2BJAWlfBcJDEIKSAWZAxboj3Qaq/bFsOyg7aAiQ3Ray20F3O1DTgGIHV1dQZigxCkkfkILgmFD2M4He8Y9ijDEfilfnr/XtCPsgpB+GLqKIMaJt20P1x/n5OXLO7/qumx9o2JjkQgg1M3sAJymlEwAnqjoTkQkRjYmo7bquK6XEy8tLO9DfgwUgxhhjjDEG//qv/8rn5+cupVSpaiMiExGZMfPcOTcfjUbTyWQyHo/HtpXsFss5I8aI3W6H9XqNzWaDnPO3qj2OB5+b95MCh/ZGzAx1CoUHtO7bXcURKCUgpr4iZAg9NOe+KsQ7ILv9VHVzG6hCRCHUV/GUlFC6iNLugLYFdx04JiBlKDsIMxwxmBSOGQIFYeijtX+esONvjDFv3T782AchzEApGCpABCIFXdeBmTAajZBSPGxwMbcKEZEjIsfMKKVMvPdTVZ2p6gzAlIjWOefdYrHYiYjz3tsL8fdgAYgxxhhjjIH3nmOMYTQaNQDGIjITkdMY40lKaZZSalTVqj5uuZwzVqsVnj9/jqurK1xfX2O73aKUvo/RceWHhR/vN9oPhFBA9xM8eHhbCng8AouAZb/r9OjvopS+nVLOQCJbBL8lhBjFOeyqCqmqkH2AiPYh124H3u3gmgZU12AiMBEcETx5FO7/e4VCgL58aP98YcffGGPeOj1qQ0iEw2szM8E5B+/dMPfDgdnBWtXefiLics51znkSY5ynlE5CCFvnXNt13a7rum2MsXvX9/M2sADEGGOMMebDRo8ePSL0bd5DjLEhonEpZaqq85zzPMY4FZFKVfn/+mbm5umHYwpyzofe0PvwY7PZIKV01FqhZ+HH+08BkOpQCQIoE0QJ5BxcVQElg4sMM0H6m5YCzRnatqAUIcmjOI8i5eWAdKBfHDc3jhJQiJDYIbJDAvVhVoxwbQu0LdB1oK4DMfftVZxD5gJWhgNBhyxMjp8v3t2PZIwxH4z+aVdf+bjPoPsAxDkP5/pT9ZQittstmqZBCGH4d9vHdNuoKpdSqpzzOOc8TSnNRWQNYJNSWgPwpRQ7sN+DBSDGGGOMMR8uevjwId+/f5+//vprD6AKITQxxomqTksp85zzLKU0yTlXImIByC2jqhARtG2Ltm1xdXWFq6srLJdLbLdbdF13CDuICCJiFSAfiMPxHRaylQhFBMQMDh4kDUgAp3Ko+EDJkBShuxpIERI7lBCQpQAKOCngfQhibiQhQiFCBvWDzXMGxwjuOmjXAW0LahqwcxDnwN7DO4YoAMah6kOBvg3W8NaqQIwx5u06Pl/rEYhoPzcC3nsQMUrpN7xcXy/BzJhOp2iaxgKQW2ioAKlKKeOc82yo0J+VUlallJH3PkynU1ZVAgAispP338ECEGOMMcaYDxM9fPiQP/vsM/f111/7EELdtu2IiMYisu81Oy+lzEop+wDErpxuGdV+MOb19TWeP3+O5XKJ1Wp1GJT5+teaDwftt45iCMrQzwIRBQQKDQEqAhUBjRJQcj8TpG6BpgFihOSMTvr/VtChyuirRexv6WZSDMPr+zBLYwScA2KEdhHoOqAdQhDn4LwHUkDwvg9Hqa8A2XeVL+i7qIHIqkCMMeYt27e/enm+1r9lZogInHNQVbRtiydPniDGhPV6g7t372KxWKCqKmuLdcuoKqtqiDFOSilTEZnFGGfOuWlKadw0TZVz9ui3KOhQ0W0vyd/BAhBjjDHGmA/Pcdsr3zRNAFA750allGlVVVNVPSGi09FodNI0zZSZm+HrzS1QSkEpBSmlQ8urJ0+e4Pr6Gl3XHSo99hfRx5UfgIUhH4xh4ZqYXw1BCBDQsF4u4NyAcoZ2HXg0gmy30KZByXn42+mHpHspULWhqzeXglXBpYBTgmMHiXEIQDpo20F3O1BTA86DfQC8h3qHygeQ23+XIUt5lz+KMcZ8gF7OACG8LOTsh6Lvh6R3XULXXaHrImKMGI/HmE6n32p3am6+YSB6XVXVpK7rec75NISwFpFrVR13XddUVRXQX6MJ+hBELAT5NgtAjDHGGGM+PIR+pxAvFgsPoGrbtmbmUUpp7L2fVlU1m06n87Ozs9lsNps2TVN5760F1i2gqsg5o21bbLdbLJdLvHjxAsvlEpvNBqUUMPPhItiCDwPgZSssAEoOAuoDEamgKUGrCmgaUNO3SNIYISkBIuCcUVKGpggUW1y5qQgAax9UlZyhnJAdQ2MHjRWkbaF1Dew6kA+gqgLXFagIIAXQ/u+iACggMIYQhOy5wxhjfiz787eXbwERhnNAKRmlCGKMKKXAOYfdboec87u8y+b3xMwuhFCPx+NpznnnnJsT0QzARFVHIlIxc/iv//ov17Yt/fznPy8A2EKQb7MAxBhjjDHmw0KPHj3CV199RX/0R3/kcs5+NBpV2+22EZGRiIzrup6en59PHzx4cHJ+fj4/OTmZnpyc1CEEqwC5BUopiDHi+fPnePbsGZbLJdbr9WHex3734N6+EuTVtgrmQ3J83AX9okph7ltZeQ8XPFBVQAjgqgKqClRVoLqG5gx4B3JsrZBuOFKFA9CUAiaCS4TOO+Q0tMPq+pu2LbiqQHUEYgJCAtU1kAuKYxQiFCiECKSCofW4McaYH8mr52sEZuqrMYnBLIeZIMz8yqYXc7uEENx0Oq3v3bs3m81mabPZbNbr9XK3201yzqOcc5NSqsbjcXDO5X//93/HEIIQYKdkxywAMcYYY4z5wHz55Zf02Wef0WazcaenpyGl1BDRCMAYwKSqqslsNpvev39/ulgspicnJ6O6rp1VgNwe+7kf+7ZXMcZD+LEPQEReNrCx8OMDd9RSAwBE+8XtwgxyDhQCEAJcXUOrul8Mr2tQStAYQT5AmaFEsAnoNxcBcKogCKgUEFFfxeMzNCZQ2/bhVn0UdoUKFCpQTAjMKACyYzgCsip430YNZM8hxhjzIzsONvrwA1B1cE4O53z7lqgxxldCEXPzee95PB5X3nvXNE0MIcxTStOu6yZd102aphmFEOqu66rdbkfL5RK/+c1v9Msvv+xfmi0EObBdfMYYY4wxHxb+8z//c/fs2TN3enpaAxiLyDSldCoiFymly9lsdrlYLC4//vjju+fn5yfz+XzivWfnHMGWN2+8nDN2ux2ePHmCJ0+eYLlcIud82AH4+i5ACz8M8Poiysv2GioKSD/jg0RAucAN70MEWgpcTvA5I8QIlzNYbDrETUREL/sfDmsiOuwcZgABgFeFA4Edg50HeQ/2vg+5iCDUdzkTEMA0hF5Hzymqr35sjDHmjTs+n9u/f7zJRVXhnEMIAU3TwHsP59wwL8SqQm4LIiLnHIcQPDOXUkq3Xq+3bdtudrvdpq7r66qqOiJKbdtCRHS73erFxYU+ePBAHz9+bCf4A6sAMcYYY4z5gDx69AgAaL1euxBCYOZaRMY552lKaSoiExEZl1IaVfUAmOwK6VZ5vTe0c/+fvXPpkeQ6zvYbcS6ZWbee7pkmh7QEXaDV0DsB2hiGvdDeK/4ezvwCL7yyVtrP1j+AhteEYAgkDEGwDcGfbiOyp7vrkpnnnIhvcTJrqmu650KRnOqZ8wCFuuWtqjJPZcYbEa9BGrK9939KESkXwIXnkKEaZPR3EGYkY8DOAXUF7WtQDKAUQX0PtBvAWoAJxGV/Olh2hE4ighVBFQNsC2iKMCGA+w5GEpQJGCp/1GUzdIaCtYIhwBAgyhAQlLKQMnbCKtGWQqFQ+PbZbWs6Ph6re8fHbdviq6++QowRXdfh3r17OD4+hjEGxpSc+FsAAVuRi1XVppSqEMIkxjhLKc1jjPOu61oAxMwqInJ0dCQPHjwo2Sg7FAGkUCgUCoVC4R3i888/p7//+7+npml4s9m4lFJtjJmq6lREZiIyTSk1McZKRKyqlhr5W8LY1irGiJQSVHWb5TdWeOze7z8uQkgBeBZQEWTPCCJCIgIZA3EOXNVAE4GUgBjBfQBt1iDnQMZAQc95gdCzhX/3H6hwLaQKowqPCFWBxgjuO1DooFCod9Cmgfgq/7bWYij6gDEEw5SFMQCGCJJ/+SJ+FAqFwnfEKH7sV3DuVoKEEPDVV19hs9mg73sQEbz3sNbCObetCikcPsM1mSOimpmnxpg5ER0x87LrutZ7ryGEtFgs4vn5eTo9PU1vepsPiSKAFAqFQqFQKLxDfPTRR/Q///M/XFWVnU6njoiqQfSYDbdpjLERES8iRou77a1AVbfZfZvN5orp+f50+xfKRfwoXGHYFxSDIToIxAw1BmLMEBivc/VHiJCuB6oqVwsYBjgLJrKzT7EqWLX0zzsgxn6GJJKFqZSASNCUoNYibWaQ9Rpa1dBBAFECYBhsDcxghm4sQZXABIgWCaRQKBS+a/bP9cY2VyklpJTQ9z36voeIoKoqWGuRUsJsNkPTNFtfkMJhw8xsrfVN08zm8/kRMx9774+JaJ1Satu2FSIK6/U63LlzJ/73f/93+VF3KAJIoVAoFAqFwrsDffDBB4TsA2cAeBFpRGQWY1yklBYiMkspNSmlKqVkRaScPN8CUkroug5Pnz7d3i4uLhBC2F4IA7jSKqEIH4Wb0MHHYVcEETYQa5FUwSpASqAQgb4H1Q3ghwoQZiRmBDZQIpAqfIo52F4qQA6H4begncf5BYKGAG07yGYDrdfQoXc8mEDWgJ2FsQZ2qC5TCIQYCQImQiq/c6FQKHwnjOd1u8/H+7ECWFWRUsJyucQf//hHtG2Li4sLnJ6e4r333sN0Oi0CyC2AmW1VVZN79+6lpmniZrMJm83mIoTQhRA6VRUAvXOu/+qrr8Lp6WlQVSKi8qeMIoAUCoVCoVAovDM8fPiQjo+P6Q9/+AM750wIwYlILSJTVZ0S0YyZJ8zcEFEFwBT/j8NmvLCNMWK9XuPs7AxPnjzB06dP0bYtYowAsL2w3RU/gOIBUrgBoq2ZtRKgTNnvwVoIkF8TBcVRAKnBVQ21DmIsoknonYeAQJJgVMApoYRXbgeaEqTvIW0LWW9AxkKshRoDOAdTVRDnoTa33RNjkAAwCKKSW2EVM/RCoVD4ThjP4/aFkF3DcxFBCAFffvklLi8vsVqtQESYz+domuZNbXrhNTDGmKZpamst13Ut6/U6nJ2dnV1cXKy6rluLSOecW8UY19PptJ3P5/zo0aNSmjlQzkELhUKhUCgU3hE++eQTrFYrPjo64sHg3A9m540xZjabzWanp6fze/fuTY+OjuqqqiyXlLCDZbyYXa/XOD8/x1dffbWt/Fiv1wghbC+G90WOfaP0QuE5iCCqUCiECYkJafABSc5DqgpSVUDTAJMJZDJBmkwRJ1PEZoreVwjOIVkHYVOC4bcFVVBKoL4DVivQ8hK6XCKtVtDNBmhboOvBMYJjhEkCI7ptc8bYGVtKJUihUCh8Z4yix+5jItq2uEopYbPZ4PLyEufn51itVogxbo3TC4cNEbG11tV13dR1Pauq6gjASUrppOu6477vFyGEiapWbdu6tm3NJ598QqWdcaZUgBQKhUKhUCi8Awwnv9T3PTvnDAAbQvAiUonIZDKZTI+Pj2fHx8fzu3fvzk5PTyfT6dQ554oAcqCMba/Oz89xdna2FT9G74/di+B9E/RC4VXR0dDcGCgrVA0SM0gEVNdAHyDNBDJbIN3ZQI1FWq+RkgAxgPo+L6MIILcCGvxAuG1hmSFMiEQQZ6HegZoaHAJMiIAXqOQqEEMEZgLGChCgiF6FQqHwhtitABnPCcfzwRjjVvgo7VBvDzSAbAdSEdEkpXTU9/1x13WXzHwRY5zWdV2JiGNm89lnn/FPf/rT8eT/nb4IKAJIoVAoFAqFwrsB/eIXv+AYI282G+O9t13XuRhjnVKaNE0zvXfv3vyHP/zh/O7du/Ojo6PJbDazRQA5XGKM2Gw2ePLkCf785z/j6dOn24vZ3cKdMbNvV/woQkjhlRkEkFEISQoQM5IIKEZwHaCzGVKIQBKo94j+EqltQZsNOCYolWHk1qAKjhFoN6CUECULGsk5aFWBNy1M34NCAELMhuk8tFkBwESQK4srY02hcBDsef1sXyvB77eK/QSY8Z6IYIyBtTkMPFaFlELvWwunlHwIYR5CuNN13ZKZnxpjpuv1urHW+hij3Ww2/PjxY8E7Ln4A2fyyUCgUCoVCofAWo6r06aefmt/97nfOOVellCYppWnbtndTSqeq+v6dO3dO7927d/q9733v+N69e7Ojo6PGe8/GmDHbqHBghBCwWq3w5z//GV9++SUuLi62F77M/Jwx5q73R6HwSmyDJ5zdsml4jbO5OYnm9kcyVBgRQcAQAEkUEAFJgk0JJJqbIw2jSRlUDpRR8ALy78iEZC2CcxDrwN6DvQM7BxgDGAbYQJghnPcB7I09hULhO2RsfYksSEIVjGdDOBPBgHaGdHo2Ho+CSBFGbjU3tT3dbYvqvUfTNFv/j90qkXLaf/iklCTGqJvNRlNKQkTRGLMSkVWMceOc64wx/Y9+9KOw2WzwT//0T/r48eN3+o+5VIAUCoVCoVAovOU8evSITk5OzNHRkb28vPTr9bomooaIJqo6UdWJiDTGmMpnbFVVJVHmwFHNrWdSSgghIMa4zfArFL5JdEgcFACDwzWIGWwNknOgqoI2EZwSNAkkBmjINwoBIYTcWgkKmxKspOF54dAYxY8IICoQRdGFgNj3oL5DajdwbQu0Ldg7iDVgY2AMw4iFNbRtfyWq22qQYopeKHwHXCt+5KZ0o9iRD0XdHqfjMU/AtlWhjMsqx+ytY0x+2a8CYWYYY7aVwiKyTaIZzyGPj49LVcgtgZnZWuvn8/kUwMJau1ytVgtVnQ0+II0xpj4/P98YY/THP/6xqKoQ0Tt78lUEkEKhUCgUCoW3nAcPHtDZ2Zk5Pz93zFw552oRmTLzFMB0qAipY4xeREwxy7sdjJUe4203a2+s9hgvcnefl8y+wuuguxnB2GmDBYDYgJ0DVxUoJUiMQN8D/QTUdUCM0BjRpYikiqiKBj1YBSW8crgkIgQ26IxBT4QEQGIEdz247yFtm1tkeQeyDmwtjDVwdhBfiaEqUMJW6CoeMIXCt4eqbis6MN6L5PMCVTCNFR+DTw/tCJV4JnzKcJ7AQxD9nY2UviVcV/kxiiAhBJydnaFtWyyXS8QY4b2Hc27bJqtwuBhjuGkaC2DaNE0/nU6P/vKXvyz6vp8vl8uZiExVdeW9X3vv5de//nX66U9/mvAOt8Iqe3WhUCgUCoXC2w2dnZ1x13W2qirftm1tjJmklGZVVc2qqpoR0fzk5GQ6m81qa601xpTY5IGyW/GxXC6xXC5zdv1e26vd2y5F/Ci8Ltt9Zsgc3gbKmCHMSM6CvQOih2lqoO+hbQtqGkjfQysPTXUWUERhFdlAXTXfMATrSkXIQaG7N5EsboUsfkjbgjYtyFcg50HWwjgL62zeL1S3vbbHZZRs8kLhG2ZMaBjHUc0SNWFoUYjchpBHwZqwnQ4JAGVhkoihBAgINNwDz+7L8Xv72K0C2RU/9v3huq5D3/dgZsznc4QQSvvCWwIRsbUWTdMwM9eqOqmqasLM05TSlIgmxpgmpVTP5/Nw7969sRPeO0sRQAqFQqFQKBTeYlQV//Iv/8IxRisi3hhT930/ZebZZDJZTCaTo8lkcnT37t3F6enppGkaVwSQwyWlhLZtcXl5ibOzM5yfn2O9XiOltL2w3RdA9n1AighS+Drk+NeYNZxbpIhhCCyitaDKAymCmhrUN0DXgfo+t8MSAUSAlNCrAJKgqrAisGOgrnAwEABWhVGBSQmaEuLQ0ky6Dtq2+VZVUOdANotgxiZYYuhQNaIAeLjf7juFQuGvY/wfJ3omIufyDTB0KzBDFaz5NYgO4giAQSTBIHzAGMhQQZrvAVHKVSAYWx+W4/e2sXuut9sGa2RMqEkpYbPZoOs6pJQgIs8tq3B4UMZ47wHAxRgrY0wDYEJEU1WdDi2Oa2NM++Mf/5gBkKrSu9oGqwgghUKhUCgUCm8xj0FxOtEAACAASURBVB49osViwU3TWBHxXdfVqjpJKc3m8/nivffeu/Pee+8dHx0dHS0Wi+lsNvPOuSKAHCgxRqzXazx58gRPnjzB2dkZ+r7fVoGMF7n7F7C7GYCFwteCsG2JwqMAQoTEDLIWMSVY50F+uNUVqK9AfZ1bYYUAiR5dTFARJFXUMYIlgUvG6cEwih9eEjgCDELbByTrkLoeWmcRhLoOaFuQ94BzgPdg53J7FWbwmG2+Y7ZcGuoUCn8lo1E1npmakypIFKwAj9V1ItAYh+cyiCN4VmmnCjCDrYVyAlmTfZ2MgYIgPLS+2zNIL0fw7WK/CmRXADHGbD3jrLXPeYYUbhUkIial5FW1TilNRGT0AakAuM1mY4Cdv+N3kCKAFAqFQqFQKLzFfP755/Szn/2MY4w2hFB1XTchoikRza21i+l0Or937950Pp830+m0cs4xF/fDg2Xs27xcLvH06VNcXFwAwLb91U0QEWToB14ofG2G3Se7gRCUAOVcCcLOQpKDqSpoVYHqGhQCeKgc0BghMUFjQpAEpIQkAlV5Ry/FDxeG5nY6kqBCCCmBYgLFCO17pLYFbTaA87kF1ugDEzzUGAgTmHMG+ZhFrpTFlOIrUCh8TfbEj5zODbBSrvRICUYUlCIoCTT0oJQr7zBU4dHoBQYAxoCsBZwFnIMYA7EKtWZbYbJd9ZXNKO2wbhO74scoiIzeccaY7fspJazXayyXSwCAGwTtcklw+KgqA2BV9apaA5gM1R9N3/d1CMFXVWV++9vf8k9+8pP0prf3TVEEkEKhUCgUCoW3mI8++ohEhLuucwC21R8A5gDm3vtp0zST2WxW13Xt3vDmFl6CqiKlhK7r0LYtNpsNvPdXejvvZ/ztvlYofBPkIHY2z01EgGGQGJCzIO/AdQ0KPShGUAiQPgyG6AmSImIMYBMhiaGl28ZhsfVlURAYSQRGBIgRiBEyCiBVDXUbGO8B74GqA1UePATMjGEkw0NlWs5S1511lABqofAa7Fd+DEblDIVRgJPAioKHMRchZD+mEKAh5raDKYEE2QSdGWAGeQ+uKyAmsPcY7UGYKIsjQ7L42AZrPHaLCHI7uMkLZDRDTyltTdHbtsXTp0+3z2ezGeq6LgLILUBVSURMjNHHGBsAExGZpJQmbds2zjkXYzS/+tWv+Fe/+tU7e+AWAaRQKBQKhULhLUVV6dGjRywiNqVUMXMjIlNVnaeU7qSU5jHGiYg4VX1nT4hvE6PQYa2FtfZKht54kSoiz4kfhcI3yjarnyAKEDOSMYCxUGfh6gok09x+RQQIATK0wSJf5QBdjAAHvOOenAfO4Ho/ZI9rCEAfkGwHbDYw1gLOg60D+6EahAyYGOwtmAYPEOZnrXTGAOqb/WCFwu1B9VkrOc2trBgAi8IqYCTBSoKLCaYPoK4Hug6y2UD7DtL1efyNCRJjPg6ZAWvBTQ3ualBdQ+uUfUMAqDHZR2Q4ryAAafQUK8LHreJlIggAhBBwdnaGruuwXC5x7949fPjhhzDGwNoSNr4FkIgYEfEiUqeUpiIyJaKJiDRd11UiYpumoc8+++ydbYNl3vQGFAqFQqFQKBS+cejhw4f87//+72axWFgiavq+PwJw7L2/671/bzKZ3L979+57x8fHJycnJ4umaSprbakAOUBUFSKCruu27QlG8/MQwnMCyL7xeaHwbUB41k6eaJQxhj70qjAYetMngYYITbntFVICDzeTEowk8FgGsuNjUzgABlPkRIQ0mJsrDbETY/KNTfYPsBZkTDaIYUZighBDmfJrw7xlZCoUXs62TRXGdlc0iB95bLUATBLYJHApwYUA2/ewXQfTteBNC6xWwGoNXa2gmw10vYFuWmjXQbsOFLP/UjZKp9xSixhkGGQMiM322AVytHR7/JZx+lax6++x+3g8XxQRxBjRti0AwHuPxWKBuq4xmGwXDpiUUur7Pq3X677rul5V+7quW2NM65xbiciKiNYhhP7k5EQ++ugj/fTTT9+5v+Mi5RUKhUKhUCi8XdDDhw/pH/7hH/jXv/612Ww21mVjj4qIGu/9bDqdLiaTycnx8fGd6XQ6G4SPkhhzoKSUtr4fFxcXuLy8RNd1UNWt+LF7IVvEj8J3wTajFEDSIcDCDLEWWnkoFBojKERQswH1HdB1QN8D1kGshViLGA2IEgwURqXUgxwYrAorApciEBkxBAgbpLaFOgc4D/hsgg7nAGsAa0Amt8ESHYRZIpgh8CYolWmFwo1s29Blr6VR+NgKIKqwqjAxwYQEmxJs38N0PUzbAW0L3bSg5QrUtqC2ze2wYoKk3P5fiQDvwZK2SjYRQNZADUOZATZZ8DAGCoWhPJFobolVjuDbx3471LGqOKWEGCP6vof3HpvNBiGEMk7fEoiIjTGuaZrJ0dHRnJnXIjIXkWkIoRGRCoBbLBYGAD948OCdrAIpAkihUCgUCoXCW8Su+GGMcXfu3KnOz8/rGOPEOTebTqeL+/fvH5+ent47Pj4+WSwW86H6ozT5PVBijFitVnjy5AnOzs5wcXGB5XKJEMKb3rTCu8xOVjAACOVWWGoZojb3jA8xG2fXFdDlG4Ue6D009Oijgw5m6D6l7Duxk/lceLMQsgDiRIAUYYjQMaM3BhICpOsB14K8B/kW5DxgGDAMdhYmWYhVQBQChTCelQ0VCoXnGce/HY+PbdsrERgVWBGYmGBDhAkRJgRw28F0HWgQP7Bpoas1pG0hgxeIxAhJudpOmaEpZtFjWxHwrEKAmEEmhwsJgJAOFWC5Emw0Ydddb5/CrWO3FZaIbFteGWNKNeYtwhjDTdO4u3fvzqqqCovFIq5Wq8vLy8unl5eXU2aumdkbY9zR0VF47733RFWViN6pw7cIIIVCoVAoFApvCapKjx8/plH8qKrKr9frWkQmIjJNKc289/Ojo6Oj+/fv31ksFkd1Xc+cc4aLy+HBMrYlODs7w1dffYWLiwuklLaZebs9nUu2XuG7ZLvvIWcUKxNEDdTltknU1JCUoHUNdB2o60EhQvseEjyQsjGvptyKxSaBKeG0g4KhcCrglDOHJTJCMEAISF0HOIe4XgPO5soPO3gLVBXUWjhnszCGZ+mmZZwqFDJjqysaDMbHtGwAMJLFD6MKEoFVgGOAjQk2BtgugLseJgRg0wKbDdB20M0GsmmhbbsVQGIISCL53AF5rDbeIw7rVMmttTirIGDiIQgOqAqsMVAGYBSqz9phEUZD9Dfz/RVej/E8kZmvnDsy81YEAXLlcdd12Gw2W8+5seK4cHgwM3vv3XCfqqqKABar1WqeUprGGCdE1CyXy4qI4g9/+EP57LPPdKgIkje9/d8VpdVBoVAoFAqFwlsCEfF//ud/mpOTEyMifjKZVCmlSdu2RzHGu8x87/j4+P3333///v379z+czWZ36rpumJmppHodLH3fY7Va4U9/+hPOz8+xWq0gItuL1vGn2xdCyk9a+NahZ/3hCTl4Rrs3VZAK0AdwSqAYgZRAMQFJsvghAsQIqym3dSkVIAdFDsgOxsgEJCIEZiQ2UMrVHjlb3Gx9A8hYkHcg60DWQofqoLF9TvECKRSwFTwY2Fa+7RqcswjMeBs8k2wIsH2A7XqYTQvbtjDrDWi9Aa0Hv4/VGrrZIG02SG2L1LaQEJD6HhojJEVAZHseoeO9AsS5+oOZwcZsj1tlysIJ5Xvi0Q8IxQ/klrHfAgu42hrLOQfvPZxz23PMUfwYTdMLhwURETOztdYaYxSAbDab1eXl5ery8vJCVS8BrLz3XdM00VorX375pf7v//6v/uhHP8K74gdSKkAKhUKhUCgU3iI+/PBDqqrKpJTc06dP6xjjZMj+mYrINMbYhBCqGGO5irlFjH4fYxYegBsFjiJ+FN4IQ1BbCBDD2TzbJcA7cF1BuwrU1KDQ58ehh/Qd0A9m2rFklh48CkCzYKUhAMZCuw5iLah1uWWOtTCVB7oO7B3IWSg8MFSBGCIIsM16V5EshpQxq/COsRWJgWc3kdzyKik4JRjN95wSTIzgPoD7HtR1oLaDbnKVB7oum5y3LdKmhXQdYtchhQCJASkJRBKSDP4dzGBrEQc/kUgEA2QDdBo8QMZzDc3VIWJNFj0MIyllQVRlO/YXbhe7yTJjRYgxBjFGnJ+fI4SAy8tLnJ6e4v79+1gsFnDOvenNLrwEVSUR4RijTynVIYSJtXZCRBMRaWKM/f/93/8lY4w+efJEkG253gmKAFIoFAqFQqHwdkAPHjygL774gi8vLw0ROWPMtv1VjHFmrZ32fd+klLyqGpSmBQeLqkKGdhV93yPGCADbTLzrpi/CR+FNohiuopkgICRSkLNAsODKA1UFqiqgrkFtNkOntgPZDmDeZhoXDhjNfh4YPEEQA7Q30MHQnowFXG5/Zdou/94+ZvHDmBx0BWCIIZyrQYYeO0MbnfL7F95udKfCbRQ9cgVI9tshEVAScBJwjOAYc/VHTOC+B/chj5tdO5idb6BtBx28P6RrIW0H6XtI10NSRIoRklKuvsKgYxJfaaXJmmOgowDCbKDGgtiAhwoQQwSwgjgvx4AgNB7H3/lXWfgr2G1DOFZsju2tYoxb8aNtWxARFosFJpPJm9rcwmswCCAmxuhjjPWYAOecmxhjmq7rOudciDHG09PTd8oQvQgghUKhUCgUCm8JX3zxBS2XS+O9t0TkiagGMI0xzlV1NviANCEELyKsquWS9UDZ7b98cXGBy8tL9H0PADDGbAUP4OqFbOmtX3gj7LTRUGYkVYAZEIF1Fsm6LIA0DdAHUN2B+h5ceWhrQcbk6Ql4R67DbyeKLIAkyeb2JgCBIV0WOECcW15Va9CmAXsPtRaGCGoMhAjGGqQx6xiAlOzxwjvEWPlEGASP0eBcJbe9SgKOKVd6xAgOAdQHmJCFD+6Hyo92g7TeAEP1h3SD90ffQ/vsz5NiREoJIgJVyecHudxqqOQwWRQRAUvamp8zEYSHKhAiEAFseBBAGGR4MEQnsGJoa/dGv9bCa7KfLLPr7TEKIJvNBgAwm83Qdd3WH6Rw2IwVICEEH0JoUkoTZp4CmAGYMnO3Xq97EYne+3h6ehrflQSqIoAUCoXX5WUj4wvff/jw4Te4KYVC4Zvmth+j4/Z/8sknePz48XY8+vjjj/XRo0fjNGMC3NsG/f73v6cPP/yQnHMmhOBjjA2AKRFNRWQKYBJjrFNKTlWLAHLA9H2Pi4sLPHnyBOfn59tMvBDClYuUIngUDoHtfjh6PAyvKZAziL0DewfxHqapwV0H9B2wzi2SyNpBRKGifxw0CkLOUocINMbsARIMtOsAa6FdC209qOvAXQfyHmmoAHFskAwjAUgYW2E9y4gvP3vhrWYIMm6rPoZ7owojCpPSIHrEXO3RDa2uhhs2LbTL4gcNBufadlkA6Tto10NDyCJITEgpQkQgKSGpQvRZpZ4SQZMBRMDjWE2chWgAAIGJYEwWPMia7ANhHWJMUEtQUkTVXCGiCkWp4rqtjAHwXW+50fdjvBVuB6pKqsopJTe0PJ4w8yylNBORmaq2VVW1McY+pdQ/efKEAaQ3vd3fBUUAKRQKN0GqikePHhEAfP755wQAH3300ZWzmt///vf005/+dPv8D3/4wwvPeh48eIA//vGP5czoG+arr746uO/0/Pz8jW3T0dHRt3oNfXJy8tZco9+/f//KZ7ltAsiXX365v5/RD37wA/zzP//zldd/+ctf6snJid6/f1//9V//VY+Pj+Xjjz/OXQCI3orfc/jtCACvVisLwBtjmkH8mKnqJKXUpJSqUQB5s1tceBExRiyXSzx58gRfffUVVqvV9mJ03/S8UHjjDAEwDG2Mtp4OlM1yjbUQ58A+t8LSugJ1Fch7wHmAxwqQgzudKeyRM9ZzxrgmhsYIMgEIBtIy2Fmg9UDbgqoKNBjpGmshxoCZYJiz38DQ/moUzoAighTeMvYyq6+YnauCRbPJeYywSXLlR9eD2w7UtuC2BTYbYJPvtd1Auy4bm3dZ9MhVHz009EAI0JSG21D5IfL8gUWURUzNniCkijQYoBPyMZqIQNbCWJvHbusgzsEahopAOPuGJFUQZwFbyxF8a9jN+t/3A9n3nIsxbm+7IknhICEiYiJyzFwbYybMPCWiuapeisiamVfGmHY6nRoANMT83vqDtwgghUIBQFaKHz16REMPQJydnfHjx4/pZz/7Gf3Xf/0X//znP6eLiwuaTCa0XC6paRo6OTnBBx98QACwXq+pbVuqqgpVVREAtG27/Vf03hMA/O53v8N8Pr92G7que6V/0dls9trzvC7f1nJvYjqd/lXzn56eXru9fd+/SRHiTa36W8F7ry96PrJara6dv6qq1zqpqKpKl8vl68zyyuu5vLzcPv7d7363fVzXtd67d2/7/OLi4rXXv7usrz3zC9gdVwDg7t271HUdjeOOc46ePHmyfey9V++9tm2r9+7dk8lkkvq+T23bpl/+8pep7/v08OHD9PDhw7eirvvLL7+k6XRqqqqyxhgHoE4pTURkoqoTALWIVKpqSwusw2ZsgXV5eYmLiwtsNhs0TQPnHKwtp/CFA2TMAh4CfOOgKsQQY6DeQYIHxwCqaqhvQVUNuFwdQq3NPiCFgyQHbRWsCoscVE0pQgOyxwfn3xl9D3R9zlb3HuzcNoOcjYG1BiIGwow4xFtk2GcU2AoihcJtJ3f0G4zOt14bQ8srUbBIFj9SylUfIcD0Aabrt+KHrlag9Trflito1+b2ViFA+x4SIzQEaAig0INjzOKHCCDDeCwKxo7ASAwBZeMRPCu+044ggwG6MCMxg70HWQs7CCBs8zitRBACzNgaC4DSUCNWPH1uBdcJGKO4MYogRIQYI1arFS4uLkBEaJoG3vtyLnqgMDMZY+xkMqkWi8U0pTQnorm1di4isxjjEkBVVZWNMZrlcsmffPLJrUuC/DqUPbZQeLchAPTw4UN8+umn/ODBA16tVtz3PVtrDQD+/e9/b+7fv8+r1cosFgsWET49PWUR4c1mw845YmZS1e3jlBIxM1lrCciDMAAYYwjIQXnv/XYjUkoEANZaxBif+yfen3Y0gt35DK/EuJ5X+mK+oZQG59zXnvd1thc3fA/jd/66vGi7X2e7ROQ7P/Nl5hcG3kXk6wbmt/MZYzSlq5WixhgFru6v+9sVQrh2nn2MMbrZbGCMuTLN2P//Jqy1N27X7jKqqtpOvz/t7jpms9nX+q5u+lzfBFVVbffBGCMxMzvnCAAPYw2rKjnnxkwm7bpOm6ZJfd/H5XIZjDF90zQdEfUxxu74+LhX1YhbXg3y+eef0/e+9z0esn4sAJ9S2pqgi8gEQCMivrTAuh2o6rZ/93gbAwtjL+ZSBVI4KHYy+scqEGVCGioAuPLQFIG6BzU1UGdjdHYebM0QkCnD0qHCABxyHx0nCQIFVJCgiAAiM9A5iGsh6zXIWcCYvF8YAzKDCGKyADL+AzGeCWZUPEEKt5ztKCZ6RTgcTc552+4q30wcWl4Nba+460Ft9vfgzQa0XILPz2EuL6BdB06CNHh3IEYghlxBEiNs6AERiCj6HW9yRT7Oso2PZAFDaWuKDmQfCA4B6LpBBCGoc4CzQOVBxmzFD1aFgYchgjXZG0RU85gAPKsKLCLIQbPv/bDbBmv0m1utVvjjH/+Itm2xWq3w3nvvYbFYFAHkQGFmruva3rlzZ8LMaTabtW3bXnRddx5CuAghXDJzvdlsPDPbo6Mj3m0b/TZT9thC4R1krPb4/PPP6fj4mAHQr371K1NVlTk6OuKUknXO2cvLS8vMZrVaWWutjTFaETF93xsiMtZaDiGYIYjGREQiwsYYGh8P96MwAhEhIqIxyCoiNP55Du9tt9MYAxHZCh7jtLvP9z/bTQH3VwnEjyWe30TQfmdZN05jrd2uaz8wftM2jMt9lWn3v8/rGMWpfV4SFP3OhaTX5IXXzbsB7l2xZF842A+Ej78lM29Fgt35Y4xXnjOz7op1IrJ9f1xXjBG6E73cfX983Pf99jEzX5n+uQ++89647pTSleUz83b9IYQr26yqyszbeZn5iqCy/3lfZTu+acb9fRxXmJlTSsYYwxg6CvBOo9oQglhrBUAE0ItIx8xrVV2nlNbWWjjn5NNPP5UnT55sWyN/W9v/bTK0KCQApus6a631yBUfjao2QzusmpkrIrLDuP2Gt7pwE+NF6H7bKwDXGqAXIaRwMIyBLzzrNw9roGKhLkGcB3kPUw3iR11vs4zBVPSPA2YUQBgKLwpVAYQQoeiZ0BqGWAc4B9lswNZChtZmai3IOhjnoTHCmCHAOpih6+CNUEaywm1lK3wMVR5Arr4wyD4fnFKu+hgrPvosXGS/nB7U9c9MzjcboGuB9Rq0vIQ9P4d7egbtewQAxlgICKzZi8fECBcj6hRBgwBC4O02DT1fsXuiK0BuZTW8RyGAjQFFAwQDdAxtW8B7wG+2IiYoD9WGGcZkf5/x+MXQUit/IUXMPHRo5/969zEzw1qLlBJWqxXatsV6vUbXdZhMJmiaBk3TvMlNL9yAMYa89/b4+LhumkZns1n79OnTxdOnTxd9389EZJJSqlXVE5E9OTl5Z866igBSKLzdEAA8fPiQHjx4QKenp/Sb3/yGHj9+TD/4wQ/4gw8+4KdPn5o7d+5wCMF67+3l5aUF4GKMDoDr+95Za20IwQ0tU6yqWmOM7brOEJExxnCMkUXEAOAh6M1DoJKJiGKMNAbDVZVGcUNVKaX0XKB8DHIOmQdjJcmVlk77gf+bgva789/EuB3jNK+SFX1Tpvj+sm7axt3A8k3r2/+MryOAvOJnuHaaFwkXr5Mx/iayy1+Wwb8bnN+ddl+sum4542sicqOQsvv6vhBARDqu57rH1y1TVbciBBFtH99U6bK73GFbr6znpm3ZXebuOnbXfdPn2ufbEkDGfV1VaRw/RMSklEyM0QzCB6eUeKieIQDCzDHmQahNKW0AXMQYPTOzqkqMMX3ve99Lv/nNb0RVb2sVyGiAzs45A8D2fe8B1AAmVVVNm6aZ1nU9vXv3bjObzSrvvXlDImXhFRlFkN1+y/viBxG9UGwvFN4Iw9Ai4z7KjMic26c4C/YOWlXgps4CSF3l9645zykcDlvvAiD3+tdcDcKJgBggvUEyLZQIhgik2WBZQIBzgLUg52C8g7UGiuwzYJihCoAJcbcdVqFw6IwZ9KMHEkZ/D+RqDx08PlJud5VNzgNMCOA+PBM/NhtQ2+WKj80a1LbQrs3vr1awlxewq2Vud8UMZz2ICEkVSAlGEnyK8CmBRXM1BikYhLDjG5YrPgiquYWVgKGiECFoYiBGUAi5HSEx1G0g1ubjlxlk7ODtxGDDsM5CjUANI9dnD2M/SmLGbWFfBNk970wpIYSAtm0B5Er8vu9fmAhXeLMQETGzqaqKjDECoGnbdkpEoxH6hIgqAL7ve/vkyRNzdnb2ThihFwGkUHh7oYcPH26vU1arFZ+dnfHx8TGfnZ0ZY4xxzpk7d+7YGKNlZrdarRwROSJyACoR8UTkuq7zRORSSs4YY1NKLoRgVdUSkSEik1LiIZhoUkqMQfgYq0CIiHJckcaKhyuCyCgW7AbzRyFhfAzgikAxvrYbZH+ZCDLyInFiyLL/2gLI/me6aTt233+V7R57cN70/nWvv0j0uW7+mwSg1xGGDqmlzr4YsPs68LyQcdM0+68NXCt6XCcU3CQejOu/TgC5bht3H++LFrvcNM9169gXQcb767bzus/wKmLBXyso7LT62R7349gSQrA74utWBBna8MFaK0QUAQQAaxFZWWu9995Ya1VVQ1VV3fn5ef/9738fn376qd5GEeThw4d0cnLC6/XaxBjt0OKqUtXaOdfUdT09OTmZ3blzZ3Z6ejo9PT2tBp+QgzleC88zVoDcVAUy3u9evBYKhwRRbo2iRFCbg3LsPbSqoH0A6hrcNOCqAnlX2qUcMmOAbHi6+0sZSXCRoNTnCEpK4BRBMQApAgSId1Dvc9VP5WGdhahmIUQVhgmi2FaDlDGtcPDsiB+MZ9UfBgAl2VZ9mJhg0nAbxA9qe3DXgbo2t7pab8DrNczlJWidfT8QAhDydGa9AnctECOUGV4EBkOFhea2Wk4SnAhIFQqFKMGA4IajdTyiFLQVQkQVSoSUgEiEGHio5hiOcGuhxkKcy9fI1gAMkGGwMzCVh6odxJVhjB8NtXfWWThs9hNsdmMIKaUrJuhlbD54xjiUUVVrrfWq2gzixyzGOCGiWkT84BXCAMZY3Vv94xYBpFB4CxlbXH3wwQem6zq+c+eOZWaTUrLL5dJMJhO7Xq9dSsnFGH0IwY1ixxAw86paD/ceQJVS8kTkRMSKiFNVhzyGjALINgApIttWNEOwkkfxY1f0wNVrqCtXvON0KaV9EeDK4yEDHLvzf10RZHx/WMULr8Bf5jNx3TbcJKy8bH37IsjurC+b/rrg/wsEit3P/9w8ryumHAovqEa4Vsy4aZqXVXZct8q8i+qN8+0G2l+w/Oce7y/3pm3eX8eLhIxxudcJIDc9ftlJ0jdxEnXDPszDsc8pJSMiRkTMKMjuehARkQzVH30IYUVEF0PFCAFIzNxWVbU+Ojrq3n//fb24uNDHjx/fqlZYqkqPHz+mL774wnjv7VDB51W1otzyajKfz2d/8zd/s/jwww8XJycns/l8Xk+nU8svO7ALb4zdDLwXiR+FwiGz23KFDSOJAQ1VAFxVoLoBNS24rkHWgYwF0TuRiPhWwaqwKYG0g8YIdB2wWQHdBrHvchusugbqGqauoV0FOAfjLCwRBAQlwPCz4GwJnhYOmkH8oCHQT6O5+Vj5kVKu+kgJHALs0KKKQ8jCx6YDtS2wGbw+lkuY5RL27CuYy0vwegkSgaYESnFbOYLBUN2MraaGg4R0x2ck12ehgsIjV+Jd2fQ8B6CAEiBKiKRoE9AyI8Xcmo4IgG0Bv7yMWAAAIABJREFUw5AhESMLIJzbYXkH0yRoEsBip7pk+E7GypjCwbNfATIytHCGtXZrij6emxZuBSQiNqVUpZQmMcapqk4A1NZan1Jy6/Xanp6ejiLIN3L9fqgUAaRQeLughw8f0qNHj/jBgwd8dnZmAdhxcAPgich3XVcNg2CNLG7UIlIZY6qqqurFYtFMJpOJc65SVT8a5lLuGW91aIUlIhZZWWZV3XqBIA+0uwLIcxUgw+Nt0Pym6osXiB/b9/arRl70Bb2sMmJXBNlf1ssqBV607t1t33v9hfO9bsXI/nv7q33J93OtALInDL2MQxFBdgP2V97Y+b2em/ZFy9mdd5j/RiFgECiem/RV5t+dd78K5boKkd3Xrptu/Az71TD738N1Is51679h+uf4Jk+edrd7Z8xgERlvJqVkiIiZmSk/oCFzXpxz0XsfiGhJRNMQAoUQJKXUWWuXm82m6vt+86c//UlDCHp6eioPHz6khw8f3oYTQHr06BE9ePDANE1jYozWe++7rquMMXXf9xPv/cRa28zn8/rk5KQ+OTmpmqaxzFz0jwNjbDUQQsDl5SXW6/WuJ892ulL9UbhNKJANdRUgCyRVmKoCRKAhgEIPXc+h8zlkvQZSyoHB0GPw24YOpxc0hMcZKIG1A4IA8Jh5LgJFgkRCBEGMhWw2SKsVtGmAqsoCmHMwyFnnvA2qmexaQKWFTuFA2Q0Uj5UfoyghQ8WHyODvkcChz+2uuj63vupymyuzXgPrDbBZ5zZX6zVouYR5+hR2dZlbYWke/SAKUhmePxM7nm1TvqNn0saO6bnuToLnZlJAQIiCXPVBARHD+YUkEA3jLhGECWSGhAxrAO9gJg3UWcAa2OG45eF+d1sKh83+ueR43T+aoY/PY4y4uLhAVVVQVVRVBe99MUQ/XIiIbFVVk+l0ehRjvOz7fpFSamKMlbXWNU1j+r43n376Kf/jP/7jW519UvbSQuHtgADQxx9/TB988AF7703TNAzALZdLH0JoANSqWvd93zBzIyITVZ2IyARAo6q1iDTe+8l8Pp+dnp7Op9NpRURen3l/mKHVjBERMwQgDa4RPMbs7J3Kjytixw0Cw5Xn1wTrr32++2f9qgLIsL6bvsvtezvB/xvP3faC2q8kTOxvw6tUT9xUmfGy2V623K857dfZlu+UVwzAf61p9gSOa9d7XQbFTZUY+9Ptiwx7J6QvrMC4bsP2t+W6+fY/0774sT/NdymA7AR7rwimOwIIj2MQMxOG0t8hQ0mttck5F1X1MsZYnZ2dBQBt13WXOlS7XV5euul0Kin33aNPPvkEQxvBg75uU1U8evSIV6sVz+dze3l56WKMnojq8ZZSagDUg8jt6ro2g09I4cAIIWC9XuPy8hJPnz7F+fk5+r6Hql7xABkp4kfhVkA0eIEAGAJoyRqI90DTQEKAzudId+5A+x4MwJhL8AqQECAAAmUB0KjCqgxCSOFg2MmCFyIIgEiMKIIYE2LXQboWtNkAdQ2qqnxjAhseDNGzD0iuAkERuAqHx7ifA1fEiHwxPHh9xAibErjvYfoA0/egtoMZ/TzWG/B6BXNxAV6vgaHVFbVtFkaWl+B2DTNUe1zH7vpv4rpWdTfBBJAKVBI0ZV8RlQSksBUjhU2u5DIGxjDgLaiuQH2A9RFkI8QwDOXqkTRu5/jVvcJ2FA6D8dxyrPagoR2riKBtW3z55ZcQEYQQcOfOHSwWiyKAHChERIPIMblz587Ce3+02Wxmy+Wy6fveq6qt69pUVcV/93d/N8bx3toqkLKXFgpvB/Txxx/Tz3/+c/bem/V6bTebjWnbtjLG1MaYWQhhCmBqjJnGGBeUTZDmqjpLKU1FpDHGTJxz88VicXT//v078/m8tta63cqOsfXMeD+8tj3H2g1Q7ogHLxM2tp/jVT/wKKIMj1/5i3oFAeTKe68igHyddb/Oe9dt1zexzm+DQxFBvqk/7Rct52UCyIvmf9mJxU2Cxyvy0ulftMwbqkhem29DABkeX6n42hVDxkFht3x7OGkXZpa+72er1crHGNcppcvlcjll5qauay8itu/7OJvNGAA9fvz44MUPABjaHdJf/vIXA8B5772IVMiid4NB4B6q/iyeCdWFA2Ss/PjTn/6Es7MznJ+fo21bpJR2vZiuzDNepBYKh8i4t26ldCIkZhhrkUQhdQ1NAokREiMIuQpAiWBDyEEWAVrOmq1VAQnAgwhSODwUhMSEji16tkjMEFGg68GbDbhpctufqgIbA2Mt1Npt30kF5Qxyyi4EReQtHArPZeIN4geLwKqCB/HD9gG8aWHaDty22btjvQFt2lzlsbyE/eovMKsVsF7lCpIYgRDAfQ9O320SNiG3sXMQcAoQSUCiPF6rIKiiI0ANQa2BGoZxDlTV4LYDVx7kXBY+mcDEMBiO4Z02WOVIPmxuSqqhHUP01WqJ//f/Ai4vL7BcLgFkY/Smab7rzS28AsxM3nu7WCym3nvtum61Wq0WzNycn5/7tm0dADudTs1vf/tb/slPfnJrWkB/HYoAUijcLrYVD48ePSIMPhuLxcKEEOx6vTZffvmlExF/cXHhnHO1MWaiqnMimhHRDMCMiI689/P5fH7knJsT0TylVFtrmzt37syOjo4Wk8nkzmQyqb33ZhQ6hnVvqzf2g2h7osTXCva/ThDnbQrivU2f5V3nmwz8v+6yXjVI8F1ldXxT69mvANl774ogsjuG7IggSkTadR0xc1vXdW2M8apqmZmttTy0zCIAePDgAR48eHBrAsvHx8d0dnZmicinlOqUUsPMk8lkMiWiaV3X0+Pj42YymXhmNrfhM72rxBjRdR0uLi62LbD2fXB2M/Nuyz5aKOx6gRDnfvLikEUQEaQ4y6boIcKECA0BaNvcmiUmBDIgFbAkiEopDjhkhiFp/HeWJJAQQH0P7TrIZgPyHlTXUGPAzoKtgeFcBcIE8GDBfCsyEQpvL2OVx/B01++DVMEiQJIsyMYE7vN+Tl0PWm+ATQtqW9B6nVtcrdfg5SX48hLm7Axmvcom6DI43yTJra6u8b/7tiEARgWsBCUBkMWLPmTRmqyBbBzUOpAxoLoCtw2o3QCVB1sDEgvjLAQ6tLPTq8fvYLheOFxuaoVFRPm/Ogn6/hKqAmMs2ra91q+xcBgQERljjPeejDGN974RkYaZm6FTQJVS8qrq1ut1+Oyzz+Tf/u3fht57bx9FACkUbg/08OFDevDgAf3iF7/gn/3sZ/z5559ba62LMXoAvm1b3/d9DaDuuq4iookxZgJgoapzZPFj1jTNwjm3ODo6Ol4sFou6rueDCXo1mUyao6Oj2XQ6nVVV5a21pU1KoVB4KyCiEEKonHPWGMPGmG3Jdl3X2nWdAsAXX3yBBw8evNFtfVU+//xzWiwWxlrrRKRq23aSUpp672eTyWR+dHS0mM1mi7t3784Wi0XtvTdDm7DCAaKqCCGg6zq0bYu+72EG49HxInRoofeGt7RQeHUUzwLZQ1gNiRnRKKx3ud98TFn0GCpBpO+gbQshRgwRURQUA0xUKA3B9bfy8vz2QwoQAUYUIgmScma7dvk31baFeA+uapCxgLW5DRYzxHBuncO0dX3ZBuR0WHCh8G2zl1wwZh1mLw4FpbQVPShGIEZQCKCuB7oO0nZbAUQ2m62/B6+WsEMFCC8vcnVI6N/Up3zGTmuvrfHSgCEC83D8GgtxgwCyXkOqCrqegJwFMcFUFQwUSS2MAdSYbQutNAbVy3F8qxgTbcYKkJTS9ty0bVuEEJC+44qlwmtBzExDwp9DNj+vjTE1gFpEaiKq27b177//fi8i8cGDB2+tolUEkELhdkAff/wxA6D/+I//MH/7t39rfvvb39qqqqoQQi0ikxhjo6qTGONkaHfVqOpURKaqugAwtsCaMPN8sVgsTk5Ojt9///2jo6OjqaqOhum2rmtfVZUtQbJCofA2QUTKzOKci8aYaIyJAJKqxr7vk/c+bTabbReO29D/9KOPPqKUEg9ieA1gklKaGWPm8/n86Pvf//7RvXv3jubz+WKxWNSTyaQIIAfMeJE53o+33ZaP1z0uFA6d3aolJYIw53YpyEbCUnlQVQF1DZlMoPMjpC5A2CK1LWLXwwK5Rz3tdpYvHBqE7IVQI8JEwDCjCz1i6KF9nytAnIdUG8C5HDy1BkR5vLMgiDLYcN5Xtg7PgxBSxr3Ct8lz4geBoYAIeGhzRSmCQgTFmKs+ug66aZG6Ftp20LYDNhvo0AKL1qtc9XF5AbNewbUbUNeBbkPgWPNnR4rQ0GcvH2tArUdar2FWK5C1ADOgAobmsRpD5d/QvlDG6g99djwXDpPrWmGN56M5eczAGAv7/9k7l+W4jitrr70z81zqBlSBAEVJ/h3Rgx7Qw576BRzRUz6PwNfoV9AD9NR+gB6aHT1xt6IVli3ZJIG6nHPysvc/yHOKRVpu32SzQOYXUQYEkyAK575XrrWsPX69cP5MMfYArKpWqtowc0NEjTGmevXqlQMQrq+vH8CJ6a+jCCCFwnlDYwkv//73vzcAzOeff272+72r67oSkVZE5imlZYxxkVJaVFW1nM/nq6qqlsaYxYkI0qpqKyLtYrGYX15eLlar1eV6vV6sVqsZETGyQszjymjzbndHoVAoPDRUVUREYozivR/6vh9EZCAib4wJRBScc9Fam4ZhkMePH8v//M//nL3wMfHkyRP65ptvjLW2EpFGRGaqOlfVRVVVi+VyudhsNrPFYtG0beustVzO7efFtKIuxojD4XCME1BVGGPeih8A8iC5iB+FB8cYgUXjRwWyCwR5ICbOwtQVMJZj62wGXSwAAInyIFwlQSODmIGHMDj8SCEABgoSyQPe6CHBAsOAZLPoIa7KMVjO5pdhsDH5BQI7k+epxFn+ODnfPZgLdOFBoargaT97p+zcQIGk4JSyAOIDEMaoq2EUO/aHHNvXv3E68TCA+wE4HGD3W/B+B9MdwN6DUgLpA1lorZLPuWNPiXoP6XtQVSHtDzDOASYLHcdBOfPxfkUB8DtD9SJmnjfvFqEDgDEGqgqRLHyICLquw263Q13XsNYeX4WzhVJKVlXr8bmxAdAYY2oAfd/35rvvvmN8oAmUZc8sFM4XevbsGT958oS/+eYbc3V1ZS8uLqwxxgGoATQxxsVYZn6pqisRubDWXiyXy83l5eVlXddLa+08xtiISD2+qqZp2svLy3a1Wi3n8/lsPp/XZSBWKBQ+REREQgih6zrfdd3hcDjsh2Hoiah3znlrrbfWBmttNMak//zP/9Sf/exnDyb79JtvvqG6rs0wDC6l1KjqbBTGF8aYedM07Xw+r5fLpTPGlPu+M0NVj70f+/0e9/f3OBwOiDECwFsPnqd/p1yyCw+RowsEYyk6EYgEgIE6B7EWVDlw20B8AGZzQDR3SKQIWJsjk8BlcHbOjMPjLIIQNCWI91DbA8ZAKwe1FqhrqHMgm4enZAzIcI7SMYQEc+yOUcUbJ0ih8EMz7rOTOyHHXQkM0dj1kfs+KEZwiNm94ce4q/0BOByg2y2074GuA/UDZBhAwwATAujQQQ57oDuAhh48XuMfBKqA5H4SxAjxHmQN1DtInyO+4Bx4On7d5AqgLIJwdvwxAGWGTMLHKI6Uc/n58m7XHBHBGHOMYg0hYLvd4ve//z0AYLlcom3bIoCcKacOkBBCLSKNqrYAmpRSbYxxTdPwYrH4YA/KsmcWCucJPXv2jH/yk58YAPbJkycOgBORWlXrvu/bGONcVZcppQsRWYvIpYis67reXF1dXf/4xz++vri4WLVtOxMRm1KyAIyIGGOMrarKLRaLuq5rWwYphULhQyXGmPb7fffy5cv77Xb7++12+/thGO699wdrbQ/A930f7+/vIzPLzc3NFIH1UOBhGAyAKoTQEtE8xriMMS689/PxBtd8X4F84f2jqvDe4/Xr1/juu+/w+vVr7HY79H1/zFQusVeFDwkd/1c4D8AiMRQErRxM7cC+gg41TBNAsxaIeaU1/AD4ATowtKRtPBhIFSYl1H6AIUJQhTcGyTrI4QCyFmpzBBYMg4wFGwsyBsZaCCmYKXfHnFQTlHNh4YeCMDosNe9gjLzfMjB2fShMElCI2bnhfRY5hgF6OIAPHWS3g97fQw8d0PfAKJCQ99AYwcOQe41iehMB9WDQ7ACRBI0RMAHqDaQfAOuQDgeoMbnvgxl6EpWkoxAyxkwcf9d6IoIUzp9pm/Ho6rHWIqWEruvw61//GtvtFq9evcLnn3+Om5sbNE1Tzs9nyLgdOaXkUkrNmCYzGxfPNdbaqmkac3l5ybe3t3R7ews8rGfiP0kRQAqFM+P29pYB8GazMcYYZ4ypUko1MzfDMLSq2lprF8aYlTHmwjm3VtV1COFyGIbL9Xq9ubq6enR1dXV9eXm5bNu2BUCqyuMAjACwMYadc8ZaWx4jC4XCB4uqJu+93263u7u7u7v7+/s7Itqp6sE51xORd86FpmlS27ZpLH57EP0fqkrPnz/n/X5vnXOVMaZl5nnbtsuLi4uLxWKxdM41RGRRAvPPiinyahgGbLdbvH79Gq9evcLd3d1R/PiDqIhC4aFzEoEyOUAAZEMHM2As1DmYpoaGABoaqPdjufAAHfrsFPEWyeTBJKmCoGWQdqZMfSAEzSIWM+IwIHYdkqvAzuX+AGvHIaoFpk6Q5GCMAUDjFUzzZi6DtcLfyuj4UOSOD0yCxxiDxZoj3FgERgQcIng8D6HvofsDqO8hhwN0vwd2O+h2CzkcRvFjFG5DgMTRARUjVNKDGyceY8BEYCRBU0KKMQs6vQWNAohw7u2BtWMnCGXxw2T3BxONrj/CMcBwdHgVzpd3XSBTDBYAeO/R9z289xARXF5eYr1eF4H6jFFVFhErInVKqQXQxhhnfd+3RFT1fW/ruv5gN14RQAqF82E60fBmszGffPKJ67qu9t63RDTz3s9EZBFjXDLzRVVVl6vVar1ara6YeR1jvPDeL5fL5cVms7larVab1Wo1a5qmea/vqlAoFN4jYwfIMAzDfrfbbbfb7X3TNLu6rg/W2t4Y41U1fvvtt+lnP/vZQ3J/HK8ZRGRjjFWTWWw2m4vLy8vL9Xp90bZtO0ZffbA3sw8NEUEIAV3XHcWPly9f4u7uDvv9HjHGY6Hk9xVRFgoPmu8RQY57uDUgV0HrlCOwmhoUWiCEvKq6qiGVRwoV4ih+mJTAmgfthTNkFKhMAkAE8XllvA4DdBiQum6MvjJQw1BngcqBqwpG5HhFVlWQ5mG1ngyvC4W/iGnfGR0IU+zVKLMdB/2cEowqOKZ8jvG57wNdB+064HAYhZA9aL+H7nbQ/R56OAA+Cx8IAYgRFBOQYu7QEHlwYu3UgWJFICKQGCGchQ71A2J3ABuTB+POgp07ukHAudvHTNFXyL97Q9nVpRjL0d/rOyz8Kd4VM5gZMUaklND3PWKMsNZiGIaje7lwfkyLoVXVikgNoFHVWUppBqAZhqE2xtjtdstPnz4lVdUPTcgqAkihcB7Q7e0tPX36lABw3/f21atXjXOuTSktRWQFYAXgAsAawKZpmqv1en392WefXdd1fUlE85RSba1tZ7PZbD6f19Za817fVaFQKLxniEiYORJRb4w5GGN21to9EXV1Xffe++CcS1dXV/Lll1/qs2fPHoL7gwDgyy+/5K7rjPfeiki1Wq1mm81m+eMf//jq5ubm+vLy8uri4mJR17Vj5g/rDvYBIyLo+x6///3v8Zvf/AZ3d3c4HA7w3gPID5ankVeFwgfHieghk4uDKK8idhacHLStgdiCxv4IahrAe0iKGESQxgFa5T1cijj7s3ZhmnZCQoAMHqnrAM6l9sQmlyg7B7gKVNews/bo7pnOhYo8LC2bu/AXc1JsDmB0j9Ex7sogOz+s5MgrjhEmRrAP4NH5ga6DHA6Q/T5HuHVdFj4m8aPv3xY/RMApCyokAnqA13QGYFXQAGBJgBA0MWIIWQgxBsIGkQjW5ON5KpNXEJQNiBmGDcAGxNkBUo7jhwufxJxZa+Gcg7X2rfvXwnlyGoGVUprFGGcAZjHGmbW29t5bAOb6+pqeP3/+wa01KAJIofD+OIoeL168MAD4q6++MtZaR0R1VVXzlNIixjh1fKyZeVPX9VVd1zer1erRer2+Xq/X1/P5fOmcq0XEEJE1xljnnOVpCWmhUCh8vCgRBWttZ4zZG2P2RLSvqupARMNsNvPz+Txut1t98eLFQ1jp8ta1o21b03WdA1Bba2fz+Xxxc3Nz+fjx481qtbqsqqqy1hp6AG/sY2Hq/bi/v8dvf/tb3N3dIcYI59zxofLd3o8ihBQ+RE73aiVCYgZXDjJGz2hM0CSgwecILO+RUszHBFHO6xcBQWAxxWHhwa2w/mjQUcxICRoCdPB5gEp5aEbGgCoHrmuYWQuECHLuKJipau4CIUJZM174s5iupeO+N7k8csl5/m8WgVHATDFPKcGGAA4BJgRwP8D0WQBJ+z1w2OfS80MH7bIIQocDqOtzP4j3MCmCx/MYpwQ7fm96gG41Qh4asgpICCIJISWkGKBMUGYoEYgJOvZ98OSuIcpxdoZzMTYzCAZKBKWTLp/iAjlb3r3/PO0DmUSQSfiIMaLrOnRdB+dyhGGOMSycCaSq1hhT13U9r+t6aYzZMfNOVWcxxoaZXQjB/OpXvzpqxfiARJAigBQK7we6vb01APjrr782bdtaEbEA3DAMDRG1wzAsmXlFRJchhI0xZlNV1aO2ba+Xy+Unl5eXj5bL5WY+n18tFouZc8697zdVKBQK5wYRCRElZvZE1APoiKgnosEY4wHEvu/lu+++09vb2wexIO3p06f06tUrfvr0qXnx4oV1zrm+72simkSQ+Wq1mi8WixkRlSePM0NVEWNE3/e4v7/HdrsFEb31IKmqEJHjn58+Fh2r8KGhQB5w8+gAUQU5B0kCqiPUB1Db5lz9EKAiSHkaDk4JIcaxoFdggJzd/37fUuH/QhVIuUw5DcOxNJmMATkHbmvoMADDABsjJEWQyfE5gjxYlWMElpY+kML3c3q9FBmFD4A0uzBIFSwKHHs+cpze9GLvwd7D+AAzDMfOD9rvcwzWfg/0Y+F534P6HuyHLH7EBJviGKMlYAWcShZB8PDOT5OwzABUBVYoO0FizML1KOkQURY2xkJ0Gt1dXFVZyHQhD8PH+x3VLHxrET8eDO+WoU8CBxFBRHA4HHB/f4+qqjCfz9G27fH+tnAWkLXWVFVVLxaLhaquvPd7EdmllKYidFfXNf/0pz+lX/7ylx9cDFYRQAqFfzC3t7f85MkTs9/vbQjBVlVVhRBqa20dQmhFZJFSmqvqEsBKRNYppbVzbj3FXn366aePN5vN5cXFxbKu66o4PQqFQuH7ISJl5sjMAzMPxpjeGDMQkbfWBlVNy+VSXrx48RCev+j29pZevXrFVVWZuq7tarVyXdc5IqpEpI4xOhExKaVyXThzpofC074P4I+vtisUPmQUgBIg4zA8OQuqchQStQHkW9AYKQNVQBJijNDoIRCIKqoUYUVgyvFypuhRrEJKQAwQb6BMIOuAwYH6ATQM4CEPoOEslAhMBMOMXCVCIAIYOQatUDhyIoDS6PpgzcN7EskCaUrHXg6KAk4xx12lBPZjfNXo5EiDh3oP6npon1/Sjf0ffQ/y4/4aAjjk72FTRH1yLqKxY8TiYQogf8BYEE8iQEwARSgzxBiotRBrwWOvDxsDVBWMcyDnQIah1sJYm50jAIRO7n9Eiqh5ZpyWoJ/ei9JYaD+Vovd9j9/+9rfo+x673Q43Nze4vr4+LuwpvH+Ymay1brFYzAHIfD6Xw+Ew7Ha77eFwmIcQ6hCCizHab7/9ll+9eqXPnz9/EIsD/1yKAFIo/AOZxA8Abj6fOxGp9/t9a4xpQwjzlNLSGLMiohUzrwBcqOplSunCWns5n8/XFxcXj66vrx+t1+tF27aNtbZkuxcKhcIJOiIi6r1PKaUAYGDmnoh6Zu6Z2VdVFVJKKYSgX3zxxeQAOWvGrijq+94YYywRuaqqqq7rKhGpVNXFGI2qUl60Uy4P58i0Xb5PAJlW0k0fi/Oj8DGgRJAxRoWtgYqFVg5S16AYwGEGijlHXyRBY0DyAyRUkJSgKeX4mjISP2+m4WnKA2gNPpef+wHsK+jw9mDZVA5ghjE5Zscg7ysAshiCN4XWhY+YcTBL774UYGS3hxEBxQhOAvIBFEIWVUMAeQ8ehQ8aPOBz5B6GLIJgdCXp+JKhB7wHh/xnTAxAinApwaWEVgROR8EFbxwUDDxsAUQVpIARzd0mSEhEwHj+ntxcMpafw1pwVQF1lePtxjgkAcDjnyOm4+9Ex3+jHM/nx7vRrMAbEURVMQwDvPfY7/fw3qOua6xWK8zn8/f5Yxfehqy1pm3b1hhDzrlojNl1XbcEMBORhpld3/fWWmt++tOfytOnT+mLL76gB9CP+WdRBJBC4R+AqhIA/Nu//Zu5v7+v5vN5lVJqjTGNqi5CCEtVXRHRpapu6rpeL5fLy6ZpLowxFzHGBTMv1uv16urq6vLy8vJisVi0zjlbhiKFQqHwNiIiIYTU933suq7f7XbdMAxdSqlj5s5aO1RVNQAIXdcl4GFMzFQVz58/px//+MfsnDP39/cVEdXMXAOoU0pVjNEB4Om6UzhPJvfH9HF6sDy9pp8+YBYHSOFDZtq7lQjCDFECjICsAzWTYyBH1UAFJAmaIjQGSEpAEsQYIRzzcuLCeaLI018RQBIQ8+AUngFr8+B5yMIHdT1M34Oq3AFiRyeIMQYChdK4enwclpYz5EfK6QIBxSg0nHR9iI4dHwoO2enBIYKHIYsg3ucYq1HgIO+hQw/ph6MLBKMQQiFkUSQEIHiYkEUUTjG7SkbXR6UJjY4CyPv83fwdIOSuFCeCRAkCRVJFHGOsEsb+D9U3Yohz0LrKUVjWQgE4TCU72ystAAAgAElEQVTpgJI5OgB5dIWUe57zYroPnV7T/ep0DysiEBEMw4C+72GtxeFwQAjhGOdaeP+M28w454y1loloCCEsrLXzlNLMe99aa2vnnGNme3d3J//xH/+h//Iv/6Ljdn/wB2YRQAqFvy90e3tLX375Jf3TP/0TA3Dr9boOIbRENN/tdouU0kpELkRkHWO8WiwWj+bz+dVnn312tV6vL2ez2SrG2BBRXdd1u16v26ZpKmMMl6W9hUKh8IeEENJut/MvX77sdyNd1x289x2AAcAgIr5pmtD3fdput/oQbuqeP39OANgYY/q+t+v12gGoiaghogZApapORAwe+CLDD5nTB8cpO/l0FV2h8NExDTFH11NiANYgqYDVQUVAKtCUc+dpHEBq3wPOQY0Bxmx5LbfGZ8xYRD32gAAEIoZQAPwAGSrwMLzpVOg6UOVgRueHEMMQQTifK6WcNz9eVEHI54xj1BVojLzKUWus2aUwFZubmGB8yJFV3QAaeqDrsuhx6MbumR7oB0ifHR7iPSiOsVgxZcdIDDAhwsYAJzn2iiTlHiJRWBUYzb0j+MD2TQZgVVFDoJKFijCWyqdRiEyjq9VaizQ6QKhpQHUPMhaM0QGCCoYJgnxcY/z6B9W4/AFxGoV1Kn6cFqJPC3tO/07hrCDguF1IVY2IuDGGv1XVJqVU13XtVquVDSHIdrvVn//85/qLX/xC8AEcmkUAKRT+ftDt7S09efLELBYL/uabb8xisajv7+9bVV30fb9S1VWMcQ1gTUQb59x1XdePl8vlo81m8+iTTz65XK1WC1W1AKwxxtR1bauqsiX2qlAoFL6fGKPsdrvw3XffHV6/fr3f7/d7Ve2Yua/ruk8peREJxpjYtq188803D+GGjp4+fUq/+c1v6PXr1+by8tL2fV8552rnXA2gFpFaRFxKyYrIh7bw8INhGtZND4vGmGPU1buU4V7ho2AcnKlqLrlmgJTA42rhXJKrQMjFwjpG1WhVAWO2/CSAFO33vHlTQC0wlCAxbzYNBgg+r8gfRRDue1BdQdm8NWAzzBDK+8qxfLmcJz8eRvFjEhgYbwrOoZoHXElAJ+KHDTEXmw8e3A9ZXOs6YL/PDpCug/Y9Ut9lt0ffQ2PM4kiMQIpZtEsCSln0qCXl3qGxWB1j3NWxc+R9/o7+ThCQe0xUc50PFFYVIZ+ooSLHCWmyNjs+6joLTXWdBRBmMJsca5cYhhVKehSvZexxKdF258mpEAK8fS976myePi8iyHkyRiVzSsmllOqUUpNSaowxdQihPhwO7vLyMn377bfy+eefy9OnTycP54O+2BYBpFD4+0DPnj1jAGa/35tvvvnGPn782MYYZ8y87LruAsBljHGdUtoYY67qur5q2/Z6s9k8fvTo0dVms1lfXFyslsvlnIimLHciImIu5o9CoVD4Y6SUxHsf7+/vh9evX3f7/b6rqqpvmmYA4Kf+jxBCats2vXr16uxv5qb4q9VqxU3TGFU93rCKSEtEjarWkwOkXCTOl3dXz33fA+I0zJviBgqFD53jPj/9NzMEgMAgqQMrYNoIiQHwNXTIBeniHGAtYHLcCmJ4b++h8H8zyVNGBVYJSXJimUYCYsyilvfHWCI9HMB1BTYWxjCEGdYYqDWQ8dwo44y0DEw/At7q+Xjj+uDJ9TFFXYnkfoqYcrl5CDAhHAUQ6jrwbg/e70G7HXA4AF0HGXrw4KHBQwYPCR5IkuP2Uu4fmsQ7KwlWBE4T3Ch8nPKh7oVZAMkCj6gggmDkjeBDQHbkjb0qNAxZXDp0oLoBOwe1BsZagAmYjmchgKfBOt4Im+/xvRa+n3fjWU8FjyJ6PDhIVU1KqY4xNiLSiEhtra2stdV2u00XFxfy7bffphcvXsiH0ElYBJBC4e/A6PxgAFNESTUMQ+29X46ixyPv/VWMcZNSelTX9WaxWFx98sknj25ubh5tNpvL9Xo9a9u2tda6MsgqFAqFP59xNX0SkRhj9CGEgZkHERmQy9A9gGitjV3XyT//8z8/iGesJ0+e0P39PccYrYg4VW1FZCYicwCtqtYppUpVTekAOX9OV82dcip+FAofDZTja6ZVwIosgiQFyChsQ0gxgEMD8gO0bqB1nVcVVxXIujxQK7fMZ8u0erxSBSQdh8ZKBEkJnFIuou77vF27HlodQMbCWAMxBuIsNBkoM1SRi5fzdynb/kNmdAXQeJ6YCs4NFCQCqwAlAaeU465CBIcADhHGe1A/dsv0Pajrwdt78P097P0d+HAA+i47y1KChACNY8+QJEBypBZUAQVYFRYKN0Zd8fjzfRSciFBMBEbuBDGiMJAcSRYj1Jijm+soglQVYAyIsljNTFBjYK2FEiNhPO/jZJl5ETXPiu8bSb3baTfFuxYx5PxRVRYRm1KqRhGktdbORKQdhqGZzWZpt9vJ9fV1+td//dc0RjE/6JNdEUAKhR8eevLkiVmv1xaAizE2qtr0fT9LKV0Ow3Dlvb9JKV2r6iMAj+q6Xs/n883Nzc3Vp59+erler+d1XbtScl4oFAp/OWOfhxJRYubIzGEUPTwRBQCRiGLTNOnu7k6/++67s7+ZG286qW1bNnli7gA0qtoCmAFoMXaAYFyMV64f58Xk5pjKIkXkLTfIaYxLcX4UPkrG4SaQB9sM5L4Ha5FEwFUF1AFUVUBdAXUNVBVQudwFwiYLKKfnvnIcnQ25oBqoIGAlkACC3PsS09iv4AeQr7IDpOvAdQUdXT5sLWysoFagRiFQRH53cz/8FaqFEyax4+TzqUeGlcA6xlyJviV8GD+6PsY4K+r6Y9QVdR34/g72/g7V61fZCTJ0Y6yTQJMc45ym3prpZ8kfc9F6fn3cTI4Qi3xTSqpIkvuaeOxr4hBAQw89TG49A1M5wJocXxgTlA3A2RHGeCOEFPHjfDk9174rggB5MVpKCSGEt/ruCufDGINlADgiaqy1jTGmNca0zrk6hBAWi0Xsus68fPmSv/jii3R7e/u+f+y/iSKAFAo/EKpKX375Jb948cLc3987Y0zddV3jnJunlOYAFsMwrEMIN977x8x8Xdf1o7Ztr9br9frm5uZis9lcrFarxWKxaMaOj4/9vqpQKBT+YohImVmMMdEYE5jZE5EXkSAiQVXjMAwphCDX19fy9ddfv+8f+U/yy1/+kn7yk59wVVWmqirb933tnGuZeTa+WgANACciVlXL9eOMUFXEGBFCwOFwwHa7Rd/3bxVKTp+/Gy9QKHxMTNEnUM2FuMxIEDCZPDyzFuQcuK5BTQ00DahvgLqG1DUkJURVUEpgkQ82iuah8iYqJ/e6JM1isEkJCB485HgctgZUVZCqAqwDVzXUOYh14HGYxs6BiUEgMGGMw+LcF1N4uEwF50A29qiCCYAoSAUEBcnYIyMKE3Mnh0kJ7APsifjBg4eOogd1PXDYgw8HmO0d7P09zPYO3HVg73Fc2Kx45/O3PgHwJuLqYz6/TI4uByCpQlVASkchiVKCiREYBqhzUOsgo5CJKh/HYh2MdRDmHGdm+ej0mX63Uw9UGZ6fB993j/purGtKCYfDAa9fv4YxBjFG1HUN59xRICm8d8gYY5xz1WKxmInIvO/7RVVVM2ZuVbWx1noR8Skl07Ytffnllw/+ICwCSKHww0DPnz83m83GtG1brVarerfbzVR1nlJaqeoyhHARQriKMV4Pw/C4bdtHTdNcPX78ePPo0aOL6+vr5eXl5Ww2m1XW2nJsFgqFwl/JKIAc3R8AJgdI8N7Htm2jMSYNwyD/9V//pS9evDj7acmzZ8/w4sULds6Zvu9dVVXVMAyzEMJCRBYYI7BEpERgnSEiAu897u/vcXd3h9evX2O73SKE3FcwPTyKyPHvnD5YFgofDUSQsdhYMA7LxygsWAM4B67zYJzrGtw00LaFBo8YQh6+QWG9z46ClN7v+ym84Z34HKuKCjkOK0WP7AfJHQBkOLt6pqL7qgIZBlsLNgaWGWoYkQmJAKU8VDt2yJTonIfJqcsDWShjKCgpSBJIcuQVJwHFCCuSHR8xD9vZZ/cHDQMwDMDgc/xS1wGHA8x+D7Pfwe63sPvdKH4M4HKe+IuZ3B81AEzl75q3T0opi9CjCwR9DxgLNQYyitgwuSSd7FiMTgTi/LnQxy0unTPvCh+nX5/uY733eP36NYgI3ntsNhtsNptjNFbh/TNGlZn5fF5vNptF27arrutWIYRlSmmeUmqJqDfGuBijqeuanj179r5/7L+ZMmQtFP526NmzZ/z06VPebreVc649HA4zVV0S0cp7vxaRyxjjJsa4CSFce+8fzWazzXw+33z66afrTz75ZLHZbGZt21rnnPnT/2ShUCgU/g8mASQwczDGeACBiAIzh67roqoma628evVKv/jiCz13S++LFy/o+vqaD4eDadvWjWV1MxGZi8hCVeeq2iDHYBlVZVUtMVhnQkoJXdfh5cuX+Pbbb3F3d4e+748CyB+jbL/Cx8rkBBEgD0OJAOajCGLqGmhaUOtBIUBTQowRqprFEkUewL3ft1H4I0yrx2sVWMmrxyFj74IKhBnJOmhVAy5HnJExYFfBWAu1BmzGHiUyEM0VMOl0dfL7fYuFv5RJ/MBY56MAicKoHPs9EOPYFRNzwXmM4CHkj8fibZ/7J/oe0mchRA8HmMMBtNvC7u5hD3tYP4BCAEnZU/4aGNMwUWGgsOCxK4URx1J6hJCFKGYoWwgzjLE5utA50PjisROEmUeBlI9xhm+5Y8s90VlyWoYuIuj7Ht999x3u7++x3W4RY0Tbtmia5n3/qIU3kHPOzufz1lprQwiXXddd3t/fLw+Hw3y32zUiUnvv+7Ztzd3dHf/85z9/8AdgEUAKhb8eur29JQC82WzMf//3f1er1apV1QWAVYzxIsa4Hp0ej6qqugawiTFeee8vFovF6urqanVzc7PcbDbtarWqOfPgTyyFQqHwPmFmYeZkrQ3W2sEYMwDwqur7vj86QF6/fi3ffPONPoQh85MnT2gYBrbWmpRSJSKNqi6YeTmbzVZN0yyXy+Xy+vp6chKWud+ZMYkg2+0Wu90OIYS38pMLhcLbHFfzEyEhCyBkLWh0f6BtQDECKUFTQgohZ/iLgCUBkt4IKNMLb2KYSj/I+yVvB4VRhSqNw1NBGhjJ7I99AWAGjMnFys6BrMkRWcaATV4xbgAkzc4SAUp84EPgpFvjrXJz5NgrowCN8WgUs+DBIYK8zwLIKHZYP4D7Adz34CF/JJ+FUfH5pd5DuwPosIM57GH6DhzC+G+WfeWvYTqXHovnNPfykCTERNDg8x/yWcwQEJgJyViwcyBjQdaAbD7GiRlsDAxT3jVGQfPBty5/wJxGk51GuoYQMAwD+r6HMQbr9RoxxrdczoX3yyhYcV3X1lprQggzIpp3XTcnohkRtapap5Sq/X5v5/M5N03z4B9WigBSKPx10LNnz/jXv/41f/rpp8YYY9u2bfq+nxljliGEi5TSJsZ4VVXV44uLi8fr9fqTqqo2qnrpvZ/VdT1brVazi4uLdjabVVVVleOxUCgUfhgUgDBzGEvPA4AgIrGu60hE6XA4yGeffSZPnz49++cqVaV///d/5//5n/8xh8PBMXMFoBGRmXNuuVgslovFYnV5ebncbDbz1WpVV1VlylD9fJjKz6ceEO89VPWYl3zaAQLgWJBeKHyUvNN/M1YR5yisUQSRysE0DRAjKAZQikjeAzECISDECEkCVgWS5NgcEVhVWCiK3fo9cxKHNY7PprB/IAZg6KE7BhkDMQZauVyG3jSgygEuD1E5JRhroKPjQ8eB9tlf2D9mTrb9kSQ5AknHng9RkCL3eoxOD/I+d3uMwgcPA2jwMF0HczjA7Hb5Y98BPgApIaWEmAQpRsgwQPsO5AdwDCApsVd/E6cF9ZSPuloFrEBMCUDucRIFIgAhghgDthZaV6DKQVwWNbmqoJO7xxiY8QQ9FaGn8Z6oHNfnwbsdddN97GnReUoJqgrvPUIIEJEiTJ8XNMaRGWaGqlbGmHoUPtoQQmutrVNKrm1bY639IB5KysC1UPgrePbsGa/Xa57P5/ZwONi7u7uqruuGiOYxxtUUeQXgkXPuk/V6/emPfvSjz2az2dpau0opOWa2dV3bxWLhqqoqK3ULhULhB2LqALHWBmOMt9Z6AJGZo3Mu9n0vy+Uy/epXv5Kx/+Ns78hVlb788kt+9eqVef36tW3b1nrvqxBCC2A+n88Xq9Xq4kc/+tHF9fX16vLycrFYLFxd10UAOSNOnR6nMQGTAHL6UFgeEAsFHEWQcSEwiJBz4Q1DrYVWNSQmYIzFQYygvod6j+QbyNj/QcBRFLFIqCWBx46RcoY8TzglYBhylwAREjFS0wDVGHtWuSx+VAG2aaCKsTcm7y+K4gQ5Z47H3TRAn6KvJAuWpApOWbCkMMZbeQ/jPdj77PYYBqDrYYYBtN/B7HZwr17C3t/Ddh0oJYgoIgGi2T0mMUCCh6ZU3F8/MFMfSAWFFYGQAkoQFQRVDFB4IqixuQOkriHOgiuX+0GqKgshdZUdYcCb17g4pHgHzot3nzGm+1nmMZpw7PswxsAY85Y4Ujg/xuhkm1JqRKQVkSbGWBtj3DAMNsbINzc3D34DFgGkUPjLmGKvzG63c5999pk7HA51VVVN3/dLY8yliFxVVfVoNpvdOOce39zcfLLZbG4uLi4eLRaLi6qqZqrKANgYQ9Za5tIGVSgUCn8LmlLSlJLEGGW/3/u+74eUUg9gGAvQvTEmAkjWWum6TgHgnPs/JvEDgBmGwRpjnPe+7vu+VdVWVecisrDWzheLxXy9XrcXFxeNtZY/lJU6DxkZi0C99+j7HrvdDsMwHCMATmMDTjl1ghQKHzVjLA7Glb9CBGYDMQJxFqgriCQghNwD0rR55XcIkDEaSyQP01gVqgqrAgGVAegZQyJZoBLJxcnWQeoabCySc6DKZhEkNNkdUDnoifhRhI8z5dQxoAqojqXZenRqsY7CR0w5+sr7XGw+DKDpNQog3PegwwF2t4PZbWFfv4bb3oMPBzCyKKYgWGOQ2AIquZS7xPD84JxGCyrytlWdRAtCZAaCh/Z5KD51fpDLzi5qmix2pQSIQJJAyRzL0On4vQvnzLS4xxhzXOQzCSFFADl7SESsqtYi0hBRk1KqATgiMjFG/uqrrx78BiwCSKHwF3B7e0tPnjwxbdu63/3ud7Wqts65mYjMiehiGIYNET2ezWY36/X68eXl5ZObm5tPrq6uHi2Xy3XbtvOqqur3/T4KhULhQ0JVkVJKh8MhbLfbsNvt9rvdbt91XZdS6oloABAmAWS9Xqevv/5av/rqq7Pu/3j+/Dk9efKEAVjvfSUijYi0KaWZiMxTSosY4wLAvK7rtm3bejabuff9cxcyKSUMw4D7+3vc3d3h1atX2G63CCH8wXDu1AVyzvtkofAP5yT2RPAmRkWdy7EoIkBM2TXQD9DgoSFAUoLECIkJevxzERVR0T7Omek8OLp3dOhh2ADGQJgBa5AqB6oroGlgxv4XFQuhUSQDjs6hsqnfP/pOt8ckgLACLJr7PURz/FFKoBDAMeWOjlHsoGHIIkg/gPoeGHrgcIDZ7+H2owCy3eZ+Dz+86RUhhrKBcgQA2ElgKSeBH5ZTcevNFyECJEpjcX0AiMEQWIlgFcBwPp5ns/z/j24+tRZQhSggTMWtd+ac3sOeOkCMMbDWHr9WhOnzRVVZRFxKqQkhzMZOkCalVDVNY0XEtG374A/FIoAUCn8BT58+pf1+b3a7XdW2bbvf75fMvAwhXIjIOqX0iJkfO+c+uby8fPL//t//+3Sz2VwtFotV0zSNMaZEDhcKhcIPjKrqMAxyf38//OY3v9lvt9u7w+FwH2Pcp5Q6a+1AREFEYkpJQgj6+PFj/eqrr4Azno/88pe/JADmyZMnLqVUqWqjqjMAsxjjIqW08N7PvPdtCMGJSHETnhFT6fm3336L7777Di9fvoT3/piLfErJRi4U/gyIoASoYYgaiHMQUSDmGCxqm1y8G2IWQYYBEgI0RiAGJCaI5DFdXhteOHc4JqDvQCpIqlBjIG0LzGageS7FttOqcSYkjKuQy/n0bHhL/CAaHR84Oj1sEnAI2c0TIsgPoCEAfQ/te1Dfg/oB8B7S9SA/AF0H7g6wu21+dYfcDRLDW/8uq8JJysP28b+57Bv/UEgVEAElAXkPFyNqP4BldPLN54DP52obc2+LSoLIOEwHIY5OwML5MsVfTf12kwAyvYq7+bwREZNSciGEJqXUppRaIqoBOO+9jTHybrd78BuwCCCFwp/BFEOy3++d974eTwoLVb1IKV2mlDbOuaumaa7run5yfX19s9lsbtbr9aPVanXRNE1rjLEl6qpQKBR+eCYHSN/34e7urnv9+vW+67q9tfZgre2MMV5Vw3w+jyKS2raV7777Tm9vb8/6KfgnP/kJzedzs91uHTPXwzC0IjJj5vlsNpsT0eLi4mI+n8/bqqocEZVrzBkhIvDeY7vd4tWrV3j9+jWAN6vjTh8UpwfDIoIUCn8cBaBEEDDEIDtAnIVWDoh1jlHxAeqz+KF1DfEeEgLIGCRjkEQQRcAgWODtSJ7C2UGah+MkCXAOctiBx64X9R6IARQjIAlJGcyUy7RRYnPeK9Owc+z0mAQQVs2uDxHwGHNlfDiWmxvvQf0A7Xto14G6HtR1+TXkr1Pw4L6H6TuY/Q62O8D0PUjSHzg7CAqjCh7lTtL8tQc/xXsg5N+1wqjApgRVgVOFCwAbg3A4ZEeP93m7Bg9EB40JwgQhQho7m97tBCmcD6f3rtM97en9rfceh8MBdV0jpYSqqo69IIWzgUTEppSaGGMbY2yJqLbWViklV9c1M/OD32BFACkU/gSqSs+fPzebzcZsNpsqxtiIyLzrulWMcS0iV8aYK+fc9WKxeHx5efnk+vr6enR+XLZtO3fOlUiSQqFQ+DuiqhJCCPv9vt9ut90wDIfFYnFg5r6u6z6lFJxzsa7r9L//+786doCc9Vzk17/+NX366acGQGWMaQA0McbZGKe4XK1Wy/V6vdhsNrO6ritrbRFAzghVRYzx2P9xOBxgjEFd12899E0PjkX8KBT+BKMDRERzLIoxSKqAq0BVAjcNNOQOEHgP6XugriHBA8GCg0HgBM8MEkBVYKEo9uwzRgQEASVA+w7cD6AhuwB43NY0xuYYY2Aoi1w0iSDMYx9BWUH+D2NyeuBt90cWPwQmSY5EiikLH/0A4wN48Dm+6tABfQ85HEDji/f7XHzuByAGsB9g+j47P4YeJsbv/zlQBM73DanCiMAhAQI4SbBQwLq8TYcBNPgcfRZOBM2U9yFDhEQEUQUxF1HzDCEiyHjeBbIIMpFSwuFwwMuXLyEiuLi4wHK5RFVVsLaMo8+FsaPYikgtIm2MsTXG1DHGyhjjRMQsFgtWVSKiB3sIlj2uUPi/oefPnxvkY6Xquq4VkUVK6UJENimlRzHGawCPq6p6/Pjx408+//zzJ5vN5nK5XC7btq2L66NQKBT+vow3YsrMyRgTjDHeGNMzc2etPTBzz8xeVeMwDNI0jfzoRz86+5u3uq4Z4/XHe99Mpedt2y6vr69XP/rRjy42m81qtVotVquVq6qqzPHOiGmV4hQF8G4B5Pd1fpSVjYXCH0dVswOEctQRmAFrAZdAUkPrXIqtIWYHSNsieQ9xFWA8gjEY1AGac+kbTIXbZUX4g0AVkAQNAToMWQTxPgtewcJoHpYayuXLOmXOj+fUs7/ofwicuD2mCCozCh88uT5izMXmIWbRo+9zz0ffg7oB6Dug64HukAvNt/eo9juYvgP7IYtiMYJihE0RXErNzxYCYFRRS4Id73mMCngUNJDiKFiPQogfQD4XozMBDAKxgI2BGUcqOjqLyvF8Ppy6mKd73em/h2HA7373O+z3e6zXa9zc3ICIcHFxUQSQM0JVOaXkJvdHSmlGRC2AmogcEdkYowHAqioPVQQpe1yh8Meh29tb2mw2xhhj27at+76fD8OwDCFcpJTWY+zVzWw2e3x1dfX46urq+tGjR1er1WrZtm1trbUfglWsUCgUzh0iUiISY0xg5oGIhlEA6a21g4h4VY3W2rTf78/e/QEA1loehsEAqKy1TUppFmOcWWvn8/l89ujRo/nV1VU7n8/rqqrYOVeuN2fE6Uq40xfwtttjigo4/TuFQuF7mGLijquBCQQGWYuUBKapITFCaw+pa0hVQasqRydZCzUWQcfV6CkP5qrx+CtH3gNBBJTy8Fv9kAfivoZ1DgGUI7DG3gDGFJk2XvCLC+TvxluDzzGy6Oj4GF+T48OOwgcPA7gfwH0PPowxV4cO6A7Qvs9un8Me7rCD221hhz4LXppjlSCl0PwhwBhdIMhC1bS9kuTuHoxiFkIA++zq0uBhmGDZQESQmKEA5OQaUFw958O7966nhecxxmMEloigaRpcX19DinB5VjAzG2NcVVVt0zSzEMIMQCMitao6770lIoN8SOt4zn9wB2ERQAqF74dub28JANd1bRaLhRuGoSGimaouQwiXzLyp6/rRcrm8Wa1Wj8fej6uLi4vVfD6f2SJpFwqFwj8MZhZjTGLmwMzeGNMD6ImoBzAYYwIRpcPhIPP5XF68eHH2N237/Z6staZpGpdSakRkJiJzADNr7Ww+nzeLxaJeLBYlZvEMmYZBp+LH9JB4ulLuNAKrCCCFwh/nKByOThAFkEgBw4A1oKoC1QHUNNC6BuoaWlW5LN05sLWIqiAVGFU4Emj2khQeACoCiEBDFj8wZAeIDgPYOVhmRDHZacAEViBR6QL5uzIOo0+jpgjZWTVFH5mUi85NCDCDhxkGmMGDu7HgfL/PAsh+B97vgUMH7Xtg7Pqw3R7usM9/L31P1FXhfPkjMWRKBFJA0+jo8j6X2A8DUFegqgJbC04JZBg8Oj6O32v6Pv/QN1P4S18k8S4AACAASURBVJjub0UEwzAgxghrLQ6HA0IIJfb1zCAiY62tZrPZTFXnRDQbhqGNMVbee1dVlXn06BEjH4IMPMybpzKgLRT+CE+fPqXf/OY3ZhgGG2OsVbUNISxjjBcxxnVVVZv5fH79+eef30zix2q1WtZ1XRXXR6FQKPzDUWZORBSZ2RPRMIkfRORVNTJzappGPvvsM33x4sX7/nn/JKvViqqqMiGECkAtIk1KaRZCaGOMtYgYVS3XmzPldEXsqQBSRI5C4a/jLcFwcoFMx5RhsHPguob4ADQNMIogVFUg5wDnsngiAqU0dopQmaI9EAh5YIo4dn+EAPQ9qKqgzoGMyVE5xkIYEOTy62mdMY2iWeGH4/R6RifiB6vmgvMksCnChAjrA2w/wHS5wJwm18d+D9ruwNt72O09cDiMXR8JnCI4eHAMIC0rxj8kCJrdICkBMUK9B7zPUVjOgawFWwsjuetJVGFGJ8gxAqu4us6CdxfwTPe90+d/bDFQ4XxwzvF8Pq8ALObz+Wo2my1fv37d7vf7ehgGR0R2u93ar7/+2nz++eeTHvngLqlFACkU/hB69uwZv3jxwsznc1vXdX04HFoiWgK4ZOar+Xx+PZvNHj969OiTm5ubx5988sn1crm8aJqmttZaIiq9H4VCofAPhIiUmScHyMDMPYBeRHoAg3MuEFGazWay3W4fxA3by5cveb1eWyKqVLVJKbUi0qaU2hBCnVKyY2ld4UxQVaSUEGNE13VvrXQ7zUX+PsoDYaHwp5lEkCkOhaYBGBskC8C57ABpaqBpQHUDblrA+9wboAoSASTlwVv+rniAz/EfHTrGX7H30L6H7vfZ6WNtfhlzFEFyFBbBYJyRosRg/WCclJxDFVAFKwDNro9j7FWM+RVidnxMfR/7Q3Z/HEbnx24H3m1h7u/Bd6/BfQeKYex8EbAKkBK4rBj/oFBRSEzQGKFDFj6k60DWQK3N53JnwdbAjAKIqsIAmHxAdCKEF94v7zo6TmNgjTFQ1beiYMs2Oy+Y2dR1TdZaU9f13Dk3DyE0wzDUAKqUkgNg67o2AASAPMRC9CKAFApvM0VfGQA2xljVdV0bY2bDMCydc5dN01w1TXN9cXHx+Pr6+ma9Xl+tVquL+Xw+N8aUY6pQKBT+wYz9H8rMyVobmNkjOz/6qqr6pmm8cy6GENIwDPqLX/wCX3zxhd7e3r7vH/3/ZD6fk4gYZnYiUo0xWE2MsUkpVarKxQFyXqSU4L3Hfr/H3d0d7u/v0fc9ROT40DdRHv4Khb+O05X8NGXDK6AWEGdBlTu6P7htc7xKCDlrfhRAaMyeB1HRPx4IpAoKEdz3wOGAZC3QNFDnoFUFNSYPTa0dS5MVwoo34xktLpC/AR27PU6FD1IFq4Ikf0RKMCmBY4QZOx3IZ/GD+h44dEDXAYcDaH8AHQ4wkwCyvYfZb8FDD0oPMl2l8JeiCgkRyQ+gvgf/f/bOpUeOI7v+5954ZFZVN9mkSEkz48F/ZuyFQQPeGDDglbUd7zVfh82vYcCwvR1uB/DO4HyAWRnWcryx9aLEJrsemRmPe/+LiKwutijNU+pqMX5Aoqqri93VrMysyDhxzqluPe08EDsgOrD3RVSrwneu+x3QTtvHwvXx7CyGMDNyzq85QObntwis44IrzjlLRF3OufPed8zcAfDGGN/3vd1utzalJD/4wQ/meq1b9Ua2ydpG44Dz83P6+OOPzV//9V+b1WrldrtdPwzDKsZ4GkK4Z6192Pf9ez/+8Y9/+M477/zw/v37752ent7x3vvm+mg0Go2boa6uFwCZiOIcf0VEo6pOOefgvU/DMAgAffTo0a0YrE3TRDlnttbOAojPOXcpJZ9ScjnnFoF1ZMQYsd1u8emnn+Lzzz/HxcUFxnFECOG1C79DMaR1fzQafwSzC6ROyoIZQgRYC+Mc4D2o70G1VJdyBkkGdC5nzqBomhvgFsE5g6cJdr1GRhFEsvOlINk6CBvAeZCxZdUxMzIRDHNZrnrTf8AtRmu8Vf1iX2zNUjbKNa4qRHCKRfCYQhEzxhEyjMA0Ie0G8Dgg7wbY3Q5utwNt1uBhBxqGcqy2idG3A9XixEsJCBE6BaRhAFkLeA/1U4ktdB7s3N5FIKoQXPWBSDuHHxXX++0O418PXdBt3Hu8EBGpqhERR0QOgFdVz8w+peROTk4yqhHrtrlAmgDSaFxBjx49ovv37/NqtbLb7dZba/txHJc559MY4xmA+865h2dnZ+++++677969e/e+976z1jpqZ/FGo9G4SZSIsrU2GGOmww4QY0wgovSjH/0o/+3f/q3U5x77YI2MMayqJudsRcTlnLuccxdj9CklJyLNAXJk5Jyx2+3wxRdf4JNPPsHLly9hjNlHAABfvehrw4dG4w9nDqBGXdGvBIgAZAzEGBhf3B+UUinSlRKjAxGQJHCMIDO14+8WQaowKYKGKmUQIfULiHPIvoM4B+o6kHPgGqMzix/MDCZqIsgfwCx67Evk946PEpVAImVlfhZwqsfUOMJMoXSzzI6PcQSGAXnYlYijcSounrGIILRdg6cJpgqVaALI24EqtEZgyRxrZxhkLajroJ2Heg/u0v7crapIqvtj+dYWEXyPedNn6uHCH1VFCAHTNMFa23pBjhARIQAsIlZVvTFmFj98ztltNpu42Wz4Jz/5ya07/JoA0mhUzs/P6eLigruuM8MweACdqi6cc6uU0imAuwDuGWPuLxaL+8vl8my1Wp0yM7cTdqPRaNwsRCTGmMTMgZknY8w4CyA558jMabvdyrNnz/SDDz64FYM1LlcLNqXkVNXnnL2IdCLiRcS1EvTjQ0QQQsBms9lHYC0WC/R9vxdCDmnuj0bjj+PwuFHU1f1MIGNAztYIlR4sUlap124CkQyNEZhC6Y3gfahP49hRLS6QXArsxRjIcoPsPVLXAd4Dnd/3BuhcuguACeBq1j/M7LgVg4Hvmnnl9sH9WfhglXoslffCpLJxjOAQSqfHWGKudFeirnQYobsdtD6OMMGE4g6R3Q407EpcVis5f3tQ7DtekBMkBuhkoYYBa8GdB/UdKIQSYZh6qC3xapYZ+UAEQYtTOhoO34fZBXLo/BARDMOAV69ewRiDnDOWyyWcc7C2TU0fC0REImJExKmqV9VeRHpm9iLiQgh2HEfz7Nmz9MEHH9wqEaTtZY3GAdM0MQBrjHGoAkhKaaWqJwBOcs4nIrJUVU9Epmgfbeai0Wg0bpK5AwSA1BL0oKqBmaMxJgJIwzDIMAzy85///DYM0uj8/Jy+/PJLHobBEJGtgse8+sbnnJsAcuTMF3yH9v/58UOaCNJo/JEcFFqXSW0tThBmsDWlByRnUC7lzKir1HWcQN0IHuxVB0jj+Dmc5JTSNyFTQB7H4izoe/CiL0KIMSBmGGORATARuBo/tRYng6isQm/n3ytmwQO1cwWoReQAicKI7EWouefDxAyaJvA0gYYdaBihwwDsBuhuVyKwdjvoOIKmEYgBGiN0moAUizurdoo03hb0QAApLpAcAsAM4xxkLPvT3CGDGKHWAMaCFGAmyOG4CrdoBvZ7zPx+aC2sv/54CAEXFxdIKWGz2eDBgwd49913cXJy0gSQ44Jqz6SbF98B6ESkm6bJ3717d0wp0enpKT19+nRvErzh1/x70fayRqPy3//93/QP//AP3Pe9cc7ZEIIXkd5au0gpLZl5xcwLAH3O2alq6/xoNBqNm0PrAFtFRHLOWVUjEQVjTDDGBADBORfPzs5SCCGfnp7Ojvmj5vz8nB49ekT/+Z//SUTEqmoBOGOMN8Z03ntvrXXVgdhmbo4MIoIxZr8d2vsPLw7n5zYajT+SgxWm89eiCjIMtRbqBdD+ajK3TrpS34PHDrAWZNpw/laiCs0CCQEyTcjjCDOO0KEUKcNaGGsB52CZIUYAJWSisnocpT9mLvRWoPXBHPR80Bx3hauuD6QqeqRUbkMszo0pFPFjmkDbLWgYIDX6Sqrzg8epCB7TCOQESgmUIpAyVG7F0Kzx50YVUIGmVDYTgcDIs5g2TtBpBMceCAHGOahJYGvAbDGfuTOuxlIi0sZVR8a8EEhEEGNEjBHr9RrTNEFVcXJygsVicdMvs3GAqlKNYHYAPBF1AHoR6YjIX15e2tVqdSvts00AaTQqH374IS4uLqjvexYRm3P2zNzFGHtjzMIY0xFRp6oegGkCSKPRaNwcqgoRkRhjijGOwzCM4ziOKaUgIrMIEne7XbLW5r/4i7+Qv/qrvzr6/o/Z0fHs2TM6PT3li4sLIyK26zrf9323XC4XDx48WNy7d6/vus5aa2/d4PP7zHyhx8yw1u7zjQ/dH9cdH+1ivdH487CPNTIGahUqerWwXKRMuNZuAhp2IOcANriF1/ANVUhOkBSRp6n0BwwDaLGAOgcyFjAWxjlkJlhDReCo52OpP0OrC4Tq7df+uvp8AG8USr72X96G8/scU4MytmIAEKk9HwojGTSLH7G4qHiKpbdjmsAhgIYBtBtgthvQbgcdBuhURA8dJ2iYoHUlP3Lp5XGSYXICHxasN94idO/kQkpQNlBi0BRBIQIhlKjCMYD7CHERbC2YCQal/FxR3F25nujbeOo4OBzrisj+sZQSYowIIcBai9PTU8QY989pHAciQiJiANgau9yhpON0AOo6PMshBHz44Ye3ysneBJBGo/LRRx/Rz372M+r7ni8vL23f9zaE0BFRb4zpmLkzxjhmNkTUej8ajUbjBlFVjTGmzWYzrNfr9WazebXb7da73W4nIpOIxJRSPD09TV3X5VevXsnTp0/xi1/84mjFD9TUiWfPnvHz58+ZiNhaa8ZxtKenp/69995bvv/++ycPHjw4ffjw4erOnTvOWmtu+kU3XmcWP4wx+9vDAshGo/FnZM5/n8flzBBViDFQDygzhAgMQHMGxqkIIF11gDCXgoh8o39F4w9EUeJzJAQgBMgwgLsO2O3A1pb31lqos3DGlGJlKkXo6WDCX6oIMrvyvm6AcJjvMV8BvvZcvfpGmfzDPmILAI4yrPJa3FWJuqquj/l+FnAurg8TE2iYYKZQys7HCVTdHTzswNst7MuXMMMO2O3KpPbs8oixRB3lVMRIERgVOMmt++NtRQGolHLzmCBgiAJsXXV/hBJX2Bc3CDsHtQaGGSIKMQei91yK3mLUjoJD8eOw/PzQqZNzRs65vWdHCBGRqpoD8aPPOS9yzotxHLucs1uv12a32/Hnn38uH3zwwU2/5N+bJoA0Ggf0fU8pJXbOMQDDzNY5Z0XEOecMMxMzQwuScxZmvhVn7es58TWK4zA95RiH5o1Go/FGZgFkvV4Pn3/++fry8vLVNE3rlNKQcw7Ouaiq2RiTX758KYvFQj/66KOjPl+rKp4+fUoXFxf04x//mFJKRlUNM9vlcunfe++9/i//8i9PHjx4sLpz585itVpZ732bVT8CqiMJIrK/yJvFj0MHyJv+XVtQ0Wj8idSVwPPqdSWCGgMBak48kKFAjODlAtgtgK4DeV/cIkSvr9RvEzLHjypUBJoyZJoA76qzZwA5B3YOcA7qHWAdYCyYDWICiBkZCiEgV/FDcCVyFLfHgeBRrBH7/WxeaV40Dtr/m/l8rlIKmvexWr9DXLkJ9nt7dV/Mhedco6+odn3MBec2plpyPoLHATyMwFBueRxBmw3MZg338gXsdgMeR2jOe2FFpfTwzHFXpHOxuuBW5qg0/gzMDhABOAOUoAAkhFJ+Pk5AX10gUwB3Eeo82GaQzTDW7oVF0bpPzffbuOoouF6EPjukD2Nh23t1lOwjsHLOXc65F5E+hNB3XdeFEJyImK7ryHtPT548aR0gjcb3AWZWY4xYa5O1NjJzEJExhLDbbreunsCvFIQaq3L99lviYOyqX7lfP3Do4LH9fSIiYwx77421lo1pAciNRuN2oarIOcs0TdNms9ldXl5uY4w7Zp6MMUFEUtd1aRxHef/99+W3v/2tPn78WM/Pz2/6pX8dBIAePnxIJycnnHM23nszDIMlItt1nVsul/7evXvdvXv3upOTE2+MocPPoMbNkHNGSgnTNGG9XmO73SKlBACvRWAdih3z141G48/IvmMHUK5dD/MEtHPgroN4D+47YLmELJeQ5QqSMzAO4JRAuVlBbgW1P6D0ScRSwr3bggzDzoKWMeV9t24fhcVskJggxiBBy2py4KADZBbTDruagOo5AUD7K7Crrw9EEFKA6opnkYMZoYP5oXr+vxJYvqOP8cOoryp8vNbzoQoWAVKCyQJOVfQIsdyOUxGYDsQP1HJz3m1BmzXMeg2728JMY/nMw/xnH3ze1a/3fSPfzV/fOCL2+54KrGTYxBAQBASNCYgJEgK0ih8UYhFBvIfxDlYUmjOMKSZoqceXguoR3LhprnfdzQLIoRjSBJDjpHaAsIgcCiALEelVtUspOQBmGAZ+9eoVPX78GEd8ff0aTQBpNA4Yx1EBaNd1OcaYVDUYYybn3CAiW2Zeq2q3Xq/JOZd2u92Ag3EbEembtvl7f+jrObRnVOHitW/Pj8/b/PgseBw8Xt3MwqpK1lrTdZ09PT3tVquVbwJIo9G4bdRzqqhqTCmNKaVxmqbJex+qYJ2MMeK9l/V6rR9++OFRd3+cn5/TkydP+NGjR3xxcWFWq5Xt+97udjsbQnCzI9E5Z733xnvfoq+OhJwzxnHEixcv8OrVK7x8+RK73a6sRj9Y6XaIqjb3R6PxLTCf5AVlpX+SDGMYMAx2Fqbz0L6HLpeQ0ztIwwAQwTADuy24rlRv3AKqUwExgoYBVhVetUyOElUHSClEV2aYnJGthbUGiQjWGCQUsUxAV24OvXKCzNOq1QZSpu2JqhxSBRMiENcIHiIoSbkFACaIln9Zfibt3SR7J8m3LYZcj7o6FD9Ua9dHcXxw7fqgWEWPWm6OYSyxRNttWZk/jsjDCIxD+f5uB7PblY6dEMB1EUCj8XWQKqwIOmQoCFodWZIzNBURBDFCp6lEF3oP6iJMl4uTaHYXEV05rnDlzmrcHIeLfA7Hu9ddIC0a9jhRVRIRk3N2ItKJSB9jXDjn+mmaegAuxmjHceSTkxN6+vTprbmYaQJIo1F59OiRXlxcaN/3OeecnHOBmUdV3TLzQkQujTF9CIGfP38e1+v1zjnXz6ICADCzzBsRCREpMx8sLLqafPu6Ae51lWN++OB3AFeiy17UqFl9JCJ7sQMAqyqrqplvRYT7vvd37tzpAMA5Z7z3tk3CNBqN2wYRCTNnY0wkomCtDcaYyMzJWptjjEJEaq0Fjtya++jRI7q4uKCHDx9y13Wm6zr7P//zP05VHQAnIk5VbT2XtxP2ERFjxGazwWeffbYXQWZXyPUVbs310Wh8u5S55TIBlueJ61p+zYbBzgOLBXS5Qr4bEbIgE8MDZdI3ZaAVsh498wQ+qcDUyXYXA3wIsDEiWwP1vjh+5qL7LBDvigjCDGFGZi49McA+Cu1QkJidIbMI8vrjXEUOhkoVQOrPUyrxayIKopL0Iyj7piiuVqkfihNvcgb+Kddn11Zgz/v17Prg2vNhFDCq+7grmorAwdMEGkqsmFbXB+12yMNQJqRDAKaplKKPY+lsyBnaOj0avwcMwKnA1N1FCUjESDntXSAaYtmvpgkUunqOTjA5AzV6dB93CFT/RxtnHQtvcoEcuj++KSK2caPsBZCU0t4BknNehBB6a6333htmZmst/fznP7/p1/t70wSQRqPy9OlT/NM//ZOISO77PuScR1XdMbMH4JxzDgCllOJut1uP47gA0B0KIESkxpgMQK6JIcUV/ccJIHunR/2QmL+efy8R0V4IUdU6ppXXhI95ExGzXC59zrk/OTk56ft+aYzp8QbnyGF01pseV1UyxrAxhp1zxjlH3KT8RqPx3TC77DIzR2YORBSMMYGZIxFlY4zEGHWz2Rz71RB99NFH9Pd///ccQjDGGGutdc45b63trLWeiJyImK8RyRs3iIgghIDtdov1eo3NZvOVi7vDlXAz7a1sNL4NympTISoT5KiTzkxIXFwg7D1otQJyBnIGpVh6JDZr6Di0SJ5bAFXnghMFaxGtnApsSjAiIOcgzGAQKEuJNosB6j3YWrAxEGNgiCCzaIHi0Ci3xeGx7xhA3Y9mFwhQhI/qAFEuBevKBGEDNWV1s3D5vtB8e9BTg0OBZe4QOfwjq3D+B/y/7GOnUCaYFSjl5vNtdc0YBShnGBUYUXDKMDGCwwQaR/A4AcMAbLdF+BhG6G4HHQZwFUcwTaAYQTUqi0IocWRN6G/8HszdL6wCp4SYBUwCygJNVQQJERQTUMU2miaY0IFiB7IJYgxAhLzvkwBei5tr3Ci1OxcAXnOBHG5tYdDxQUTsvbcnJyeLlNLKGHNqjDlR1dU0TYsYY+ecs6vVine7nfnNb36Tgas0yWOmCSCNRuVv/uZvdLVaCYCUc04AgqoOxhhLRMY5xyklZeaQc+5DCH3O2c+OC6CsRjbG5Or6EGOMMLMYY0Tr2f1QBLmuFRy6PA5X+IrIXL5ORLS/P4sg1f3BB6+FRYRFZBY9LIC9CALAW2u79Xq98t4vRMTX53LOmQHsb+vvmH/WLLKY+THnnF0sFvbu3bsdEVnv/bf4LjUajcZrlEW+QCKiOG8AMhFla61cXl7O594bfaHfhKrin//5n2mz2fDJyYlhZrvZbDwRzeKHJyKHch5vfaFHxmzvjzEixoiU0msF6Pti3IPIq3bB12h8S8zHGsoHhMyPEYOshTgH6TpIyqCUoDECwwDtLgFj9/0NjeOmTJwCXgRCAGlZTW5VwTSA1pe176IKYarQFKG+A6wBGYNcz9HCXKOrGDK7P2ZRgkrnB2vtF6AaYzXfVvcIjCkCBzPYWqgxUGuK8GHK75AqiqPen3/+XMKO/XXh1Sr2w08KnaOzvo7q7JjvA4CZo7ZUQTlXMUjAkkvJeRaYXGKvzD7yaizOj90OWgUQ3ZWNhh14HGFDAMUAjgkktShdchGf2udb43dx6HxCOb5mcQ4ply1GaAiQaQJP3VUZeoilE8RZGBSnFRuuggphnmppe+HNcl3cmMe/1+OvWg/I8WGM4b7v/b1795bGmKnv+2Ecx5MQwnKapoUxxhORW6/XNsaYPv/8cz4/P6fz8/OjP+yaANJoVB4/fqzPnj2T58+f5+12G7uuY2utERHSojIIMydm3qaUOmttJyJOROjAlaHOuczMGVcCiDKzAhARATPvnSDGGIjIa0LHmx4/dH+ICM3fP3BocP2aiYhm8UJEjIgYACbnbGcHCBHZEIK/uLjoQgj+iy++8ABMtbrZeRMRWyNXjIjYQ0FljmNZrVbdvXv3emstW2u55dI3Go3viuqymx0gEUAkomSMSd77TETys5/9TH71q18d9YDsyZMn9OjRIxrHkZfLpck5uxBC55zrnHOdMcYDcKpq0cSPo+NNF3WH3R+zQNLcH43Gd8csOMp83HGZnC4CiEBriS6mAO260hdB1M6wtwQCYFE6AOb3zKiCcy4dFOs1KCUgJUAyIBmU7kD8BDYGsBYwxflBVZAo06e4coJUx0dd5gbClRNkX5pez/VCBGIDa4uzRK0FrIGxFrnGrwmX36tEJbaHsHePlLgsKSIIVUEEuOoLqb/vm0SQ12z7RODakcCqRfhIRfSgmErBeSxRQhwjbEqgqcZejSNoLAXntNtBtrviAhkn8LCDHQd0NWpsdnzQHKclufzeRuMPgBT7/Qg5g2oPiFYRpDhAAjAG8BSBPgLBwWhxfzAUbEztAiHMsyhtscnNQvW89ibnRxsHHy/WWq49wbRcLvN2uw1ffPHFyeXl5Wq73fY5505VvapaZjaLxYIeP35Mjx8/pmPu2wSaANJo7CEi/PKXv9RPP/1Uzs7O4iwudF2n0zRla21m5skY0zOzzznvV+POYoW1du7+kPn+LICoqhpjalQs708Mh0JHznl//zDuqr6+2R1C83NnQWS+nV8LEc1CiEFxcxgiMiJijDGGiGzO2W42GxdjtHVl8Sx8uJSSA7C/rUKPE5H5eR6Azzn7aZoWAJZ3795V730yxvTWWsPMpsVhNRqNbxmtAkgiomiMicaYBCDnnGW5XMonn3yCx48f6zGvSnn8+DH+4z/+g7qu4xcvXjjnnFfVTkR6AD0zd80Bctwc5hofih/zY/MF4HUhpNFofAsc9DgcOkHUGIhVqFeoCDR20L4DlgvocgFdLaHTWI7RnMtkXDtejxJC7RCAFo0A+8zgEnc1jkAurQDF2UOlLN06cBU/yJgigFAVPoj3Zcqqc0yVVncI7Z0euQofqOJFKUFngA1gDdg6wFqQL7dsDNQ5qLFQJ1DDUJG9K0SNQqjeV4Fy+XmHZewHGcoof6a+9n+xF0VUwUSAyH5lPeVcY6pS6fgIERwjzBTAYYKdJphpLNFWNWoIVQTRYYAZJ8g4ltX34wAbJrgQYHOCyaV/hWqvyRw712j8sVAV7pDTlQgyCyHTtBdDyNpZgwSzK/v6/ENmx22LWLpRDmOvDl3QTQg5boiInXOWmZmIegCLi4uLpaouUkq9MaYTEWettScnJyaEYH7zm9/kv/u7v3utJusYaQJIo3GFfvTRR3OcCn7605/qMAxirU3jOAZjzOic26DER5kY4+ysoFmUKDqEaNd1IiJqjFFrrVprVUQUAKy1X3tCSCl95RNg/tnz90sVSbl/XQw5vBURZmaur2+OtzL1MQPAhBDMOI5WRGwVdNx8W1Xd/SYi3cHXfZ2Y65h55Zw7ubi4SMx8IiJpuVz2Xdd1TQBpNBrfIpxSWk3T9IMQQp9S+kFKaT2O41pENgC2z58/3+Wcw7/927+lf/mXf7np1/u1/Ou//isBMABs7frwRNQtl8tTEbnDzPeMMXdTSmcxxtOcc3fTr7lxxeEF3pu+dyh6HF4ANhqNb5Ea/bMvrmYu/Q3WQhTIIqA+wYQeulxCFo0JgwAAIABJREFUT08hZ2fIKQFEoGEAUiyT6Y3jY+53+brv1Sgm3aCICTlBtxuwdVBjAC6RVzAMUgLTVf/H7PjYiw9Uys0TFyEDtT9EZxGESqwVVWcJOVd6ZpwHvCuCiC/3NTnAOYgViGEoG4gqMikyVzcIqnNpLlOvEVmz82TvPpknfEsu1z4Ci0VBWroVWKrzIybwNIGnAJ4CaBphhhG828FtNrC7LeywA8VYJphDuFp5H0Mpo45FOLExwMUIW39+o/Gno1dRbSrleI1X4oeMI4z3pQx9nICu2wsgVCOwDHOJ0mK6OpYbR8fhGPgwBqtxPNQ5RmOMMSLix3HsiahPKS1CCIuaTuAWi4UFYO/evWs+//xzfvbsmapqPub3swkgjcYB5+fncn5+jvfff18//vhjmaYpv//++2G5XE4isrPWWhExKSU2xnDOmY25Snzy3uswDKgiiKaUtGaB62Kx+J2fw7O4MTNN02tnD2stVBXjONJqtXrt++M4kjFmjtCinPP8NdevmZlZRLjv+7kvxAAwzGxV1YUQnDHG5Zw9EXkR6YjIq2qnqv28IllVFyKyFJGl934nIrsXL15MIjKmlMI777xzZq017vof1Gg0Gn8mVNXknFchhFWM8UciAlVFzhlvun+sg7HrE+PzZDkRwRgD5xy6rtt3Scx/U+N4OCx5PBRCDvs/WtFjo3EDHJz3i426rOIXWIgKNHelD2S5hN49g8QEVoIQl4njGsfSuKWIglKErtdAKCvGZ8eHqeICQMX1obX4/OAcfui8SGxAziF1PaTrkJwr+9eB+KHMIOtAzoP6Duw7kPfgroN2EUgd0Ak0Z6j3EMMQIxAxYGNgwMhQCJm9+yTXF7CP38LrMVyz6wWKUviuc9G5gkVgRYr7I6YSYTVOoFpkbtZr2M0G/ssv4F69hNttgZShOYFFoTmV/T8nQBSSUj0uSnl66/po/LkoYqaC5/2q7mfICRoDNHlImMDRQ6cRNHmQLR0+bC0oC2AEbE1xPhEhH4zL2vjr5jj8/z90Rh9el7X353ipqTicc/a1/7hLKXXGGJ9SciEE23WdOTs7Y++9PHnyZDbeHiVNAGk0rnF+fi4A5hKf/P7779Onn36afvzjH/NisaDNZsPb7Zb6vidjDNbr9f7sbYzRhw8fKgB89tlnuHfvngLY3/6hLJdLAMCXX3752syd9x4xxtdK1MdxpPfeew+vXr2inDPW6zV1XUfee2Jm6rqOQgjsnKMYI3ddxyklVlXTdZ0hIptScjlnZ4xxKaVOVeeoq46IupRSX90fCxFZ5ZyXRLRMKa02m82WiLbMvOv7PnrvAzMv52L2+bb2lLC1lo0xpjjrjnRmstFoHD3zQHq+v899PxA+jn1g/SaBRlX3Qsf1199OmcfFdQfIdcGjdX80GjfH/nMABCEtXQvMpQDbWpiug/Y9ZLWCxIRUo300hvJv51X0qi0O69ZRosygEygnKHHRxGo0DtWIqXJerudrOlg9TgeryI2BOg/tA6TvIdYVFwnqzzIGbGzp+PAeGnqoD+CuA0KAiT0QU9k6D4kJVMvYYQzgLMiUr8XKvjidAMi8op0IysUdooefJVriwCBS3B9SS85T3nd8lP6OAbQbSp/HMIDWG9DlK9CrV6CXL0HbzZXwJ7n8/0jeiywqc8RVi7pq/PmZHV2zCwSSgZwhKUFiRA4BXEvRaZwAV6PmkgXlGoGlKOJmjYIT1aseqMZ3zuG4+HAsPEfDTtOE7XaLvu/3i76MMWghIkcFiQjHGF2M0YcQOmut77rOG2McAJtSMnfu3GFrLT1+/Bjn5+c3/Zq/liaANBpv5npe/GvLv6oSuufahMYxfMoSAJyfnxMAPHr0iM7Ozuj999+nxWJBn3/+OXddR6vViruu42EYzMuXL23XdRaAZWZnjPExRicifpomD6DLOXci0tdtmXNepJSWOeflZrM5UdW1MWa9XC5H59xWRFY1Xsse3Drvve373q9WK09EpgkgjUbjT+VNg+xZCLkNXBdrZidIzvmNJdqN4+T6x1nr/Wg0bpj9JHbtcuAyqC8TzQbiHLTvoSkhpwyaJuSYQOMIqavoEQI4p7bi/bZRRSsSAVJ644T99ceUCBmEPBeT12dkw0gxI4sip4xsbY2/KgIIVyGDjAV1PTQkqA+QEMCTL7d9XyOmPMhZcI3TgrMgZwE2YGdLTJs1pbNmjsWqXSMqtY+E9v4PkAKoQt0+8ipnUI2sonECTRNouwN2O2A3ALsddL2GbDaQ7Ray2yHvdtXdoaXIvO3vje8YgoJRRAsVgeQETgkSAyh65DAB4wTTTYD3UGeh0YE7KbFvKJFxe9HuliyEels4HCOLCMZxxMXFxf49Oj09Rd/3TQA5IlSVRIRTSjal5Gf3R+0C9icnJxaA7bqOjTH09OnTo57XawJIo/FHQETH/imqAFBFHKoqrD569IgePnxIp6enWoUQ7bpO1uu1/L//9//yMAypCiFxu90GlHOErY4Qp6oupeQBeCKaY7F6Ve2Zeamqq+12e/rll19+utvt7lprT0SkizH2IYRlzrkHsFgul6t33313ZYyh5XLZqkIajcYfzKHIMbOPrTjiyKvrHL7m2bUClAuDOe4q57wXQubnNo6TN4kd7QK80bhZDo/BDAAEEJfc+OwcyDtQ14FXK+QQkFOCpghihiUA6zUwCcwtEdQbfzwCQmTGxBaRGbkKaMIEIULMghQCJOerLo65JN1aGGOhMQFdhIbSWaDeg6cOGCdQNwDOl1J0VzpDYAzIO1jnoNaWrhBrgSqGwFpIFViUGUIAiFE9omXit4o8XAvPESJ4CqUMfiyl5rrbQnYDdBiAYYRsN5ChCH3JWljfoYsBVMW+2zGKanxfOCwwhwogJS5Ocu0CCRMwWYgdIN6BnEWuIrZED+o8uEbBMWp3D9AcIDfM9Wuy2SU9jiNEBMMw4NWrV9jtdvjhD38IZv5KLHzjZhERzjmbnLPNObucc1cj8r2IeGaehmEwwzDwhx9+eNMv9xtpAkij8f1Hz8/Poap48uQJ8AYh5OHDh/L8+XNerVbinMvDMBhVTd77/ckuhGABGGutzTk7EXH1hDcrwX0IYamqyxcvXpw6505V9STnvIwxLlNKJyGEFTOfnJ2d3XHOxZOTEwWQnHNWVYmIuKRisWHmfcl7o9FofBOHkUPXBdXbMPF86PA4FEJUFcYYLBYLrFYrLBYLWGvbyqgjQESQUkKMEdvtFtvtFiEE5Gt9AYeRbI1G44Y4iDJSoKzsp7LKP1sD03lIypAs0OUSiBG5TgRrjKAYoSJlQfy1CKB9B0Pj+wFVF0jdEvNVGToAyrn0FOQEmWOpZidISlBjQCYWMcIFsC1ODxo9yPsitjkHuCJqqDEgawDnSsG690DfAV0P9aUwHfX5ykUEkVrgvhdAZqdSKqvlESJomoDdDlQFDx1HpGEATQE6jtBxBI0DZBxBOSNr6U2QGgHWaHyXzB0gFlp6cESQqwCiVdTTECDWwloHmUbQ6EqXTgjQVPpqSBVMxRW1j9S6BdcB33euj4Xn+7vdDrvdDjlndF2H+/fvt/HykaGqVDdOKdmcs5tj8q21PqXkrLW273vDzPzs2bP50DvKg64JII3G24FW5V1RejjmExIBoGfPntHp6an83//9Hy8WC+q6Lq3Xa2ZmnqaJRYRVlVEEEJ6myRhjLBFZEXHGGFcLkXoR6dfr9aqKHytVXaWUTlJKd2KMp9baOymlcbFYhJOTkxxjXBpjvKoaY4zvus4tl0tnrbVNAGk0Gr+L6/0KswiSc741Fz3XY69EBCICZkbXdVgulzg7O8OdO3fgvYcx5oZfcSPnjGEYsNls8OrVK7x8+RLjOO6dOiLylV6Q27AvNhrfV1RLwbWUL0oMFjPEGqRswV2HLAIKPTQG5LAChQCdAhAmWBFkAJpziRrS4ghh1P6FxvcHLZOxcx/BDOUMQi4xOwBSjcsCEYgZxLyPw7IxwloDYgNTXRxkXYm9snNcFpcILGOg1gC+g3YdsFoBqxW060GzCOJ96RcxDDVm3wkyr5RnEVCsgl2IRfzYbEDrdYm4GkdISkghQmMEpgkyjuAYgBhBtefm6DMOGt9LCAqjgIVCVCAqUMnImSEpAcxALTzPZoTxDuxLITov+iJ+iIBVoQowAVmq80DkeGdj3wLm8e9hN+MsgMQYEUKAtRa73Q4ppa8sJGrcLPXalHLORkRs3ZyIeFX1zOwA2BCCWa/XfHp6etTzd00AaTTePvQwcgWA/vrXv6bHjx8DgDx79oy891TL1Omzzz6j1WpF4zhyLX4nAFxPgjxNk3XOWQDOe+9DCL0xZpNz3jDzSlVXzrkVEW0A3BGR7TRN24uLiw0zr+v3+pRSd3Jysrp3797qwYMHJycnJ4R2TdloNP4Ibktp+GGM13XxI+cM7z1OT09x//593Lt3Dw8ePMDdu3fhvb/hV94IIeDly5f45JNP8OLFC1xeXmIcR6SU9s+ZRawmfDQaR0B1gVAtxiUmiDISM8haZK9gyUDnga6D9B3Q95BFjzytYLQOS1PpVbA5wQPwbbXq9wpShYWgz4BTKS6P+r35VgAkEAKVLYPK5CwRLAE+EXoiGAKYijBSStJLhBWYQYb3/SHgIoaI95DFEvnsDDLdBZYnoK64Rtj7Eoc1CyZEkOpImkU5xFi2EEGbDfjVS5iLF5DtBnmakIlBUv5GDQE0FQHE5wQXI3yOcJJhVJoHpPGdwijiR68CFgKojoUll7i5lKDMpcvGGOSxOKmo62BiKLFvORdBUAUEKqLH4firiuCNm+HQrU9EYGYYY17bmsP9+KjiB+ecWUSMiDiUOHyvqj7n7ADYGKMZhoE//vhjOuYo6iaANBpvMQddJnNMFn3wwQd48uTJ/oz16NEjAoDf/va39I//+I8AgOfPn/Onn35Kp6enZIwxp6enbIyxIQRXT4Z9Smmbc16o6hLAEsAJgMuc82lK6eTly5en4zjeYeZVznmVUlq98847d3POd/u+V2vtkpmViAwzExG1T8RGo/Eahyvs3zTJfMwTz4eZ9Ifb3PcRY8RiscDJyQnee+89PHjwAGdnZ+i6Dta24dtNE2PEZrPBZ599hi+++ALr9RrOOTDz/v25XmrfaDRuHpnPvQByXa3PqkiqIPWgvgdCgAxFANHFEhTSPuZKxwFGAQeAVWFJYdrx/b2BAFgVMBSa6Y2rxjOKAMJ1DBLBgGQQCI4UXhUdFBYlVgoobiMAB6IHVRcH1x4RAN6DlqvSIRIScBL24gd7B63iB/YOEACiwFzynjM0VBFks4Z5eQHzxXNgHJBCQLIdwIwIlLisGGGqAOJzhNeygp7b/tz4jiGUiUlG6f/IIpgkQzNDOO9jC5WoCogGbC3scgGdAkyMoJTLsSAKMnQVgQUUAbzt1zfGofBxuM1jZmbel6KP44jdbgfnXBNFjgAiImMMd13n+r73y+WyWywWnfe+q53APqXkttutffDgAcUYj1P5qLQr6EajsedQEPl9/42q8rNnz/jdd9/l3/72t/b+/fs25zy+evVqtNYOxphtSmmhqlsAGxQRZHV5eXlyeXl5mnM+EZETEbkDYOy6Lt25c4estZmZ1XvfAXAt8qXRaFznUDiYvz58/DbEDh2Wns/28JTS3kngvcfdu3dx7949nJ6e3uRLbRyQc8Y0TViv13j16hW22y2WyyX6vgdwu/bBRuNtY9/pwAQBIRsGqS358d6VEmrvoV0H7XroIkJz3pfyWhGQZAgztDlAvlfM3S7fJAIIEQwIokXMKG0cBKIyueJV4FTg8HqE1ozWKLY5PkvnlbLOQ1MurhERYJpArsRmsXMgOztIau9IdYBAtYgfKZcekhRB2y345UuYVxegcQLljORi6REhAiSDcy5OppzgJcNBW59N40bYH3cAhLQcU6JQEuSUSvxg7eXR6tpj7yHTBFedT0ZqDBaKLgjgSrhu+/XRcF0EMcZAVRFCwOXl5b4A/eTkBN775nq/YZiZvPe8Wq382dlZT0QLZu6NMV3OubPWOgD29PSUvfe8WCyaANJoNL7X6K9//Wt5/PixDsOg//Vf/yWr1UqIKItIiDE6Ito55zY55wURLay1C2PMSkROrLWnAE6rALLbbrfDZ599NsYY78cY49nZ2dlyuSTTFJBGo3HA11lrDy9yjv2C500T5IciyOwGORR5GsfFbOFn5tfcSIcCSBNBGo0jQ7UIIAdl6GAFWbufWNO9EFI28g4SbC2hZgjNEUY3/cc0vmvKRK3CAzCq8HPDgAIGJcrnmy5aSn8IIxAjESNXVwizAaUMu93CxAi+vATZEo9FxpQeBGKA67wu0ZUAUqOwNEtxo0wBPA6gcSyxbaLoiGCJIbUXAZJhRPaOl0bjKJij3WoXiAgh5wzhIoBkJlB04DABMYBiKP08OcOI7oUToJ2ej5VZ+Jjv55xxeXmJlBIuLy9x//59/OhHP8LZ2VkTQG4Y5xytViv3wx/+cHnnzp2T7XZ7Oo7jYhiGbhxHB8Baa03O2QzDwD/5yU9u+iV/I00AaTQafxLVNaKPHz+mX/3qV/ro0SO5uLjI3vtkjAnGGENEBoCz1noR6Yiot9YuVPUEwAkRnYrIRlWn3W435pynlNIEQGrvyGul7RWu0VhtbNNovKW86fC/Ptl87BPPh5Pls/gBANbar0ysN46L2b7/JhFk5tCV1N7HRuM4mB0gghpNpAoYBqAwzkJq6TR3HdB1wDRBvQd5Dw21NNokaN4HrDTeIuaV6q7GXOmBeDB/j/FNe0bpDYnEiMzINQbLgGBFgN0OPOzguMgSbPiqw4ap7Lw0/7a6QKKuoFeZHSECpAhKESoCowDFCEtzrNeVcMLQVrrYuFnoKm5O6lZ0kLkUnZCzIFNCSgRKCRQjOCVwTjCSqwBYekBI6xE4H4RHfi3wtjD34s0deQD2hejb7Rbr9Rq73Q4hBJydneHk5OSGX3HDGMN939t33nmHVqvVcrfbLV+9erVQ1W6aJlc7QWyMkfu+p08++YT+/d//va4KOD6aANJoNP4szEJI/VLOz8/zo0eP6OHDh/T8+XMOIfDdu3dtdYR4Ve2NMdsQwkZVt6q6TSkNwzBs1+v1RlV3zrm4Wq2yiIwxxpOcsyMix8yu73vrnHPW2uYMaTTeUr6u7PzYRY/rHDo8jDH7PNy7d+/i5ORk3y3ROB6uix/GmNc6ad70/EajcRwc5pGL6lWuPAC44vagrgNCAPU9KMZSwhsjdJoA54AUgcRN/3hLmUWOPyekWiJ8coSVupr9K+hX7v0uGW7+Hms+0impxtvOLEhnAJEICbQXQYA6ToaW83WNjGVVZBGI1AVEVdpW0Xpwauv+ODKux8POY+mUEsZxxDAMSCnBWothGJBzvumX/NZTI7CMc850Xdd57/uUUrder7ucszfGuJSSdc6ZFy9e8HK5vOmX/I00AaTRaHwb6Pn5uQKg8/NzevTokYYQdL1e609/+lMZhkEASM5ZjDEphJCIKBBRZOZRVXfTNI2bzWb64osvttvt9h4z3w0hrJxzy77vV++8887q9PSUmwDSaDS+rmvhWC963vR65/vee6xWK5ydneGdd97B/fv39yJI43iYL9pm8eO6CNIEj0bjyJlXHM8xdQAyMZQN2DqYrivF0vOWEyRFUAjgnEEpgGPtU2i8XfyJYwuCwqqgU8CKQiBlP4TCqMLWyV3oN/fLtD2v8X1BUISPSIyJCIEMMjOUCWTKYhOp4y5hBh1upt5ScX0QUz2eCi2G9Di4vkhtdoOo6n78/KZOx8aNU/yG5fgjImIisqrqAHgisiklKyLGGENffvnlUX80NQGk0Wh8m+j5+bmqKj158kQB6Pvvv68AtOs6efnypTBzMsYkAFMIIajqQES7nPPu8vJyl1JaA7gH4N40TWer1eru3bt3z6y18N4ba62Zo7DqB+tRn3Qbjcafn3nQfD1m6JgdIdfL2+f4K+cc7t69ix/+8Id45513cHp6ir7vYW0bst00h+/T3M8y5xgfRmC9KQarCSKNxpGhuhcvhOZYIQUZhloL7TsgZyBGIAQgRZgYoSGAYgQFD5gA5dIFQtd/dqPxNRAAg+L2UJoDtIoAMhewU7NqNN4iivuDMBFjmqPhmAFj9kIHG4Yyg40BjAFbU+4T7Z9zJUjrlcj9NYukGt89qlpELKkdLfX9OhxLzwuM2mKi40NVCQCLiAXgiMipqjPGmGmajKqy9/6o37R2Nd1oNL515ngsVdWnT5/qxcWFeu/VGCMppbxardIwDIGZo6qOzDxM0zTGGKfNZrMTkU3OeRtjHO7cuTPlnNNqtULXdQQAXdc555xtRemNxtvF4eD4uqBwG7i+2mm+MOj7HmdnZzg7O8NyudxHLTVulpQSQgiYpgkvX77Ebrfb2/Ovd4Ac7pvtAq7ROEIOMuehCjBBpa4uthbwRQCZs+b3bpBpAoUAxIAcA3KKSCLgurWjvfG7KAJIKVJ/k1jW9qHG2wdBiJCJkZiRjLmKJmQGs4EaC7UW1rkSQ2gs2FoYa4sQwkUIUaKrzhxg7/Br3DyH0Vfz7WGk7KGLuo2djxJSVUb5CLMAnIg4EXHMbJxz/Pz5c3r8+DHOz89v+KW+mSaANBqN74wqhEiNx9JHjx7J//7v/8put0sPHz4MOeegqmPf90NKaRSRMec8pJTmbRrHcby8vJw+//zzKCJxGIZwdnZ2eufOnSUzm/Zh2Wi8HRyWh79J8Pi6x4+B686U+XZeETVHK1lrm/PjiAgh4NWrV3j+/DlevnyJi4sL7Ha7vX1/voCbxar5fW2fS43GcaKzC6R2gRABxAZq62dL9tAugRaLvRBCiwUQAjRGpJwxiUAAuBhhU4SRb44tajRm0aN9MjQaBSVAqwiiXJweYAMypkZgGai1IO8hXQd4D+o6OO9hnAcZAzADZnaCMIB6HkervjkWDsfFh4vADkWPtujr6CERsarqVNUTkcs5W++9SSlx13X09OnTo/14a1fVjUbju2aOxdInT57Io0eP8sXFBX/66afcdV28d+9eGMcxAIgikogoGmOiMSZaa7OIhN1uFz7++OM4DEPa7XbJGIOu64xzznH5xGxxWI3G95RZ2BAR5JxfExGux18ds+X9UPQ4jFaav9dWPx0fswDyySef4MWLF9hsNhCRvXX/8AKuiR+NxvFzuAoVREAtRFdmqHPQnKHeAweF6BhH0GIBSQlJBCoZWctKfpJcXCCHx/2RfgY1Go3GjXE9KhQE5Vn8MCBji/hRI6/IOZC10FkA6Tpw38M4D3bzc0scVilPP4jF1RIt187EN8/XXacdih/NPX3UkKqyqhoRcQCcqlpjjBERTikdvXLVBJBGo3EjzLFYKCKFnJ+fE4DsvZfVapVVNeechYiyqmYAkZljznkchmHa7XZBVZOq5pOTE/Leg4io6zpvrXXNDdJofP9Q1X0M0TAM2Gw22O12SCntvz/fzoLCsQogwOuv902CSOO4yDljmias12us12vsdjt471/LLQaa86PRuE0cHqcKFAHE1MJd56BdhsYI6jsgRvBiUXpBUkLKGZISJCWYlMCSQbXAmuukW6PRaDS+igKQ6vpIbJDYQIyBGgOyVdSoG/sO5BzQd9CuAxYLcN+Dug7Gd2Dvi0BSI7DmXqbjvQJovEn4eFMcVuN4UNU5Amt2gDgRcTlna4wxzEzOOZqm6aZf6tfSBJBGo3HTKADMsVi//OUvFYAQkZ6cnGguJCKaVHUEsAshDDHGsbo/8pdffgljjOSc9e7du6fL5XLlnGNqn5qNxvcKEdmvwn/58iVevXqFy8tLTNO072J40+TzMYog11/TLHrM25ue07hZDsvPZ/fRN5U1tvLzRuOWoApBWZGjTFBlCCmyNYA1IO9AsQP6BAoBlDNUBJoSJAQgeESXgJQgRuAkw4rAtHN4o9FovBEBITEjssFkDIKxyMaWfg9b+j3IOhjnAO+g3kO7DrRcAqsVaLkELRegrgOcg5oifghREVZw0A14w39r43Vm58fcfQhcxf824ePooVqCbgF4IrI1EsvknJsDpNFoNP4A9Be/+IWcn5/rD37wAx2GQQHk09PTMAzDjog2KaWN937LzKOq5t1ulz/55JO83W7TdrtVVYW11llrHYCjPwk3Go3fHxHBMAz48ssv/z97b7LkRpJdf597fYrAlAOZZFGq/tokM8kksrVqszarhax60SuZtnyeAl9BO70C+QDa1gPov1Nz0TJrdbdV10CykpmJKQZ3v98iIsAgCsmhyKoEMv1HC2IKIB2IQMDDj99z8N133+H8/BxVVb1mH9Wxy9Uf/WqPTQusXW53AutqD631Oveju+yTxI9EYo9obVKAdlZyZ8GhFNgYRBugQgBCaKyw2nB0qSpIUSAYg8oYhGARRYAaqQokkUgk3kAkQs0KhTYolUatFILSEN0KINYAxgLWgKwFXAZkGWiQNwLIaAgMciDPEK1FVBpQCpGb0PMm4qnJdwLwA9utxM9PPwC9f19HssHaedYh6CJiiMgQkWZmFWNkZial1E5vtCSAJBKJXUOm06lMp1MAkOPj4wCgHg6HVQihNMZUIlLHGEVEqKqqeHZ2FqqqCgCQ5zmMMRCRYK3NjTFGKcVIYkgisffEGFHXNZbL5br6I8a4dQB61+l37jftrxK7STcrbZvwsVlxlE7aEok9o38sBppA3RgbD3pjEHwAuQDOc0iMQFVD7AriHKSq4L2HeA/2AToESEjHgEQiccMhes3qCq09lbS2V7UxqLSF16YJOW/zPhrR41XYOZwFuQyUZ20FSFMFEvIc0dqmAsQ04kcE1kvqUe8Wb+sbb1pipXOinWQdgh5jtCEEa4zRbS4Ir1arne78JAEkkUjsJNPpNAKQhw8fytHRUfzVr34V/u7v/s5/9913Yq1FjFF773UIgVarFcUYYa1VL168YGaalHjCAAAgAElEQVQm730cj8dhNBqNiMju2+BoIpHYTpcDUtc1qqpad5SB7R3rXe08b+Z/bFZ/7Gq7bzrd/taJH32v4m77pZO2RGJP6X13BYAwI7JCVBFkNCRYIMsgPoDyCigyxOWqsWwxBlFrBGaAFYT81b6XRCKRuGI68aNmRmDVHh8JwgpRa1TaIBjbVHpo3dhdGdMTPlrxI8uaxWWQPAOGg+YyywDnELVGJIYXIIisq/iANtcp9cl2hv4koW2h6F2ful8JktgNugwQEVEiYgCYzgJLKaW01iwidHh4uLMbLgkgiURil5EnT57Ehw8f4vT0VD755BOZTCbVfD5XWZbNV6uVjjGSMYa895jP5/ztt9/KcrkM8/nc37t3L1prjdZaA1BX/WYSicSHsy0w701+sftw0tMfPAeQAtB3lP6+txl83qcvYqWTt0RiD2lnLQsIaEUQ1gZiBbG1v+I6ayxZrIUYA3QzmLUGfN0EiqQY3kQiccMJRKiURtlmfIhiQDdWV1E32R5kLZQxTZi5tYBza9EDzq6FDmQO0TnELEPMHMRaRGsQdCOudFUfMcb2GJ7YNTbFj3524+b5XOpD7xydALIOQUejKawzQLTW9Ic//GFnN1wSQBKJxK4jT548iQ8ePKCnT5/il7/8pbfWlufn50pENDMTAFZKoaoqajMBhIgkyzLK89yKiDjncq21ZmYmolQOkkjsIZtVEm8SPXY5S6MTPLZ1/ne1zTcV7/264mixWKAoitcC0PvbcHPbpRO3RGIP6b63RAA1M4mJCYEZ3NqzcGt7JbYdmCsKwDZh6FFX8K2XvY8CJQB1WSDp+J5IJK4jPasroVY8JiBSE3JeaYPaWHitIVoDWoOMfVXtYV0jgjgHagUPyvNG/HAZJGuqQYI1iNZAXNYKHxpBK0TmNvy8qQCR3sSidNTdTbadyxERYozw3mM2myHPczAzjDGw1kKpNJ/1KiEiUkpp55wbDod5CGEgIlmbBaIAsLWWf/3rX0NEiIh27uuXBJBEIrEPrHNBqqoKL1++rIfD4QoAQghRay1VVQVmjkVRhKqqPDNHay201rquaz8cDg9Go9HQWmvTj2cisd90s/CZea8tozaDz/sZIPv4fq4bIrLOnJnNZjg9PcXFxQWqqoKIvGa9tml9lao/Eon9pZ8FQkyIisGiEERAIpAQwC6DdLOSnQPVNVDViJWBrw2qECAxQkdAxwiVjumJROKaIgACCJ4ZgRoxQogRmeGVQqkNausQTFMpx841YrJ1YGvBWQZ2DirLQM424kf2SviIrqn2EKMhpq340BqxEz9UK4BQa1+4w5OgEq+zuZ1CCFgul3j+/DlijKiqCkdHRxiNRsjz/IpamQAAImKttR4MBoMQwthaO6/relCWpSvLUouIqqqKnz17xo8ePaL2XGinvohJAEkkEntDK4KEr7/+Gp999pkAADPHEIJYayMRCTMLACnLEs+fP6eiKHg2m/m7d+9GY4wyxigkO6xEYi/pWxABADOv7aK2DTj3Mxl2kW6mUyd89N9L/zJxNcQYUdc1zs/P8e233+L09BTz+RxlWb5mU7ZtH9vVfS6RSLwDnaiJVgQhRlQARMAAEEJT8eEcqLVqQdXcjmWJ2njEEOFjhPMAi4C7KpBEIpG4ZggIgRgVK1Ss4JWCkGqECa0RjEXQBrGtoKPW6oqcA+d5I4BkGbgVPGiQr8UPaS2xommqR4JSryyvmBHaSpNIbfh5qvrYO/rnO3VdI4SAqqpwcXGBi4sLiAistUkAuWKUUmyttZPJZJRlWbVarVbz+Xx4cXHhVquVJiJlrWXnHN+/f38nPUCTAJJIJPYJmU6nmE6n4c9//rP88pe/xGw2EyIia61UVQVjjIiIVFUldV3TcrlUbU4I53lumZmcc6K1VskOK5HYPzYzQPr0O9C7HkbdFzw27+9Ig+hXS78C5OzsDOfn51itVuvH+9tnV/ezRCLxI+lVdkVqf3uUQgAArQFrweuQ3lciiDiHEAJiCIBEsKCp/hBAQUBIdliJROIa0LO9CtxaXSmNUplGANEa0l5G3Vld2eayrfjgLGsEkLwRQCjLIM4Cg7zN97DN5brqQyEqhcAEj+bY3FlfJfFj/2FmeO9RVRWWyyXqugYR4fbt2/DeX3XzbjxExMYYMLNTSg2Yeei9zxaLhQWg67rWxhg1m8344cOHhCYzZKeqQJIAkkgk9g2ZTqcCQB4/fiyz2UyYGVpr0VqL9z6GEGJd17JarZiINBGpLMt0lmUOAI/HYxkMBpnW2iilkgCSSOwh20L0NjM1+o/vGpv5EYndo6vQ6U7ElsslWqH9tUqkXa4ySiQSP551iC4RpPWYJwDQqvWub2Yzc56DqhpwFaSqEL0Hag+EAFIBHCMggMQAJQAjVYMkEon9prO9Cqxa8UOh1gZeW9Q98QPGNMKHbqs/WourLuScBjloMGjE5Db3I2YO0RhEaxG1hleMqBV8a3fliRCA14SPCDTZTalPvdd0GSBFUUBEkOc5yrJECOGqm3bjoQbFzIqZLRG55XJpmdkA0FprFWNUw+GQnz59yvfv3//hTL8rJgkgiURiX5GnT58KgDCZTGoAGI1G4pwLq9XKi0iw1sJ7r4ui4GfPnqEoCpnP5/XJycmtO3fuHI9GI1ZKpeNgIrFndIPN/QyQN1WD7CKb/sS73t6bSj9vpr9cJngkMSSRuEasv8vN4FrrvdoG+LY+9nkGtPkf5D1Q15DaA94jeI8qCkSagUILwMUATsf7RCKx58RW/CiUQaU1KmUQjEZQTch5X/joLK84a6s+shxqkIMHOdRg0AofDjFzEGcRjEE0uskUUU3Vh2dCJEJoxY6AVyJ1BIBU/bG3dJPC+guA17L2EruFiFCMkWKMSkR0CMG2Yeh6OByqwWDAABjNV3VnSAN/iURib2kzQeJwOPSLxQIiIlrryMxRKUVaayMimfdeX1xc8Gq1IhFhImLnnCUiEhHWWrduWMkOK5HYZfph012nePPxzlZql+2v+qzDdtt2b7PFSlwNfXFt86Ssu77Ndi2RSFwTRCDdd7q9jAQQM0ip1s8+A3LfiB++BsoSVNeIdQ1yAVEAD4BBYBFYiRAhUBqqSyQS+wxRE0BuLYK2iMYiKgWyBqybsHKYJr8D1oI766ssgxrkoEETdB7zHMjzxvqqzfoI1iBwW+nB7YJG6JCu+qPLy8MOBg0kfhT9vnY/7zH1rXcWEhEVY9Tee6OUMgB0VVXKOccAqF2AHfmaJgEkkUjsM9KKIAAgWutYlmUcDodRKcVEZJRSWVsFQt57UkppY4zOsiwDwCLCeZ5bY4zWOh0SE4ld57JZQv3A810XPjbbd5kIsuvv46bRz57Zt4qjRCLx/vS/1SICJoIwELnJAxFjgMwBvhFApK5BZWODRVUNCRESBSIRHCNMVJCYfMwTicQ1gAhgBTEWYjPAOrBphA9pLQLJOYh1INcuXdB5lgF5BskySJ4BbfZHbCs/olLwwCsBBGgFkKairhM9umN0moCy/2xmPF422S2xG4gIiQjHGFWMUYuIISINQA8GA31xcaEWi0X46quvZDqdxm687oqbnQSQRCKx/3SVIP/zP/9Dv/rVr7yI0HK5LK21SwAXALSIMAAuy9Kcnp6aGKNZLBZy584dnJycjMfjMWmt1RW/lUQi8SPYFka9DwPSmzZY3X2J3WLzRGxbFUjabonE9aMvqFMb+CsAhBof+mg0xFpIHiAhAN4DVQ2uPWIdQCFCYiN+IEZI8AComQ+ZDhmJRGKfoUYIZmuhBzmQ5SBjmmOitaDMQaxtxA7n1otYC3EO4kxz21lEqyFaIShe5y0FAsJrWR9NRV6/8gNI4sd1ob8NL+tzJ3aHtn+0rgAhIiMiNsZorbXaWqu01jwej3fK2iAJIIlE4jog0+kU0+k0nJ6eyvHxMUIIJTMvmFnHGElrDSKKRVGoEIKazWa6KArEGNkYw+2PKmmtmYiYmdOvbCKxA4jIOhCvLEuUZYm6ri8NPe9ud3ZY+9Bh7t5jygTZXTZFj83Ko0Qicf0RAJEaAaOrAIlRwCKIIYBDANUBUnuw90CMTUVfDKDggZpfWWolEonEvkEEUCNSoK3o0MMhaDQGZ3krfGSt8OEaoSPLgMwhtsIIjEG0TZVI1AriDKJuqj6i1mvxY211RdSIHyB0I6nyWpPSMfW6sFkFsnmZ2B1EhAB0GSAmxmiZ2SqlbFEUdrFYVM45n+d5uH//PomI7MI2TAJIIpG4Lsh0OhUAmE6nmEwmVV3XyjmnlFJUliWMMbJarexyuTQxRgdAG2PccDjUzEwiwsPh0BhjwMypGiSR2AFijKjrGkVRYD6fYzaboSgKhPAqU22b7dU+DUr3q1b6S2I36G+LbZ33fjZNIpG4Xqy/132/eeZGDNEaUQRRpKn2CBFU1eBqAKlqwDeiiPgaUlWAUgATJKRjRSKR2D+EGKI1YC0ky0GDIXg0hAyHMIMhpBVFmgoPB8kzhLbKg9t8j9jmJzWCByNqhcCMyIxABOFG6BBII36IoPmXCueuK9smGW2bcJTYLUSERUSFEEwIwWqtbYzRtoKIttay1ppPTk7io0ePdqL2NQkgiUTiuiEA4nA49HmelyJC8/m8+wEVpZRRSum6rl0IQZ+dnRmlFC2Xy3j79u149+7d0Xg8dskOK5HYDbz3KIoCz58/x+npKc7OzrBcLlGW5aV2V/tS/ZGEjv0gzT5LJBKCV0meIGpFEEIUIAqAEBrBY+CB2oNrv7bForoCVRWoKkHEvRdKJBKJPUKpJrdjNEYcjRGHI9B4AjUYAvmgCTFvKz4kyxCchcoyBNtYY0WtGuFD8SvRgwGPRvgIeD3fI0qT+QHagZHTxE9G32pyMwg9WWDtJq39FYUQtPfexhhtXdcuyzJX17XNskyvVitVVRWPx+Od2XgpVSaRSFw3ZDqdyjfffBOyLKuJqHDOLfI8nzHzeZZlL7XWp1mWvYgxvpjNZi+++uqr77/++uuX33333Wy5XFbe+53yKkwkbjIxRhRFgbOzM7x48QLPnz/HfD5HXdc/EDn2tXpiW+VH6ujvHpsz0baFoScSiWsK0dq+qskBoSYHRCt4rRt7l6wd/Mtz0HAAygeN/711IGsApZMFViKR2G2I2oBzhigF0bpdTFPVMRwiTA4QD48hx7eAg0PwwQF4PAaNx+DJGDQZA6MhaDyCtBUiYZBDBjliWxUSnEVtFGqtEbSC50YUWQeeE0HQtGXPuvWJ92Qz/yPZX+0+bfU7xxhVCMHEGG2M0YUQXFEUrigKU1WVms1m/Mc//pG++OKLq24ygFQBkkgkrifSBqP7zz//PP7hD38Q5xxCCBJjNM45HUIw3nu1Wq1UURQEgLMsM1VVjWKM2VW/gUQi0dDlfyyXS1xcXOD8/BzGGGitodTrhVqbgbW7zGW2V/so4Fx3NmefdcGMiUTi5iHUTEVu8kCAoBgQhRgNQgigzDX5HyGAag+ua8RVAWgLaAViQioBSSQSu4y04kfUprHuU6oRRQYDxPEB5PgWZHIAjMagweBVwHnmIK6p/AjWQJxFsBZeawStERTBE6EGIAQEkUbwkNbiSpqgcxHBa6pHOmReey6zv9q0wkrsBl0FSJsBor33jpldCCGLMbq6rq3WWud5zqPRaGc2XhJAEonEtaUVQeL9+/f9bDarAZTGmGWM0RKRiTEqAIaZDTNnWuuhUqoCkCpAEokdoxM3usHnzRlB+yYabOZK9IWPfXsv15W35X1sy55JJBI3gNaOJTZXQUwITOtg9CYAOAOqGihLUOZAhQVpDaSIuUQiseOIUghZjjAYQjIHsq4RQbIcMhoBBweQ4RgyGIDyHMib3I+gDaKz8EYjGIOgNbxiBCZEEng0x80AtPaB8sr2qieCJG4m/eqPbkn97d1FRLi1wDJt9ocDYJnZAjCz2UwdHBxQnuf05MmTbvbHlW7IJIAkEonrjEynU0yn0ziZTPxwOKxijCsiUt57VkopZrZEZLXWA2YeE9FKRKoQgicipparfiOJxE2lP/teKfVaOfRmh7gbmN71TnJf6IgxIsa4vr0v7+Gms0/VRolE4uMiIs1saHQiCIGZGrsYoxuv+xDBtQeKApxlIGsBYwCtm4FEia9mOKfjfSKR+FB6Fn2XrNC71q+u6Oz92uczIVqHOBzCHxwiDoagPAcZC2QONBgCgwGQ55AsRxzkEOcQrUUwGt5oeKUQlELQCkExPAERgtCKHkK0FpHXwgeS+HHTeVPlR+pr7xYiQgAoxqhijCaEYGOMFoCr69q1QehqtVrx8+fP6eTkZCc2YBJAEonEdUcAxE8//TS8fPmyHgwGxXw+Z+ccFUWhlVJOa50x81BERkVRnK1Wq4yZtTHGGWO0UiodKxOJK6Qveiil3mhB1BcRdplt2SX924ndYNuJVxKoEokbDr0aPmzyQIBI3Ab7KijnGlGjrkF5BspeLdE5xLoCiYBCAEk39JdIJBI/nk5QiGiyMwRo8zzaS1B7U8AxgqTtz2iFqDREaRAzRCtIliOMx5CjY8TRCJLlYOcAZ0FZ3oSct5VukuWI1iJag1oxvFYI3AofTIhM8KCmbZ34EePa6qp/LE3cTLrzvC7b8bIg9MRu0VlghRA0ACMiLsboRMR67421VpVlyXme78wGTIN6ievEznyxrojUb7iEL774Qp48eRLKsiStdaW1JmaWrgJEa+2899l8PnfffPPNsCgKTCaTeHR0dDAcDkdJAEkkrpZ+9sKm+EFE6wqKfRuY3hQ99qntN4nLTrw2rcsSicTNohtgjFGgWs982HYAMkYgy8B5Dsoz8GAAKUYIVQ0mgvAcqijAwYPCVb+TRCKx7wgAD0JNjECM2AszBzeXDAJDYOoaWiKIGWEwRMwHCM6BrQWMbkSN4RBxMgFGI8A5RGMBZwHrELtKN2ObYHRrETTDK27CzIkQiBCJEUBNXhLwutjR9Z+I0iDGDac/eW3TBitlgOwmrfjBIrKuAAkhOO991uaBGCJS1loOIVD7nCvfjmlQL7G5B+7lkWU6neL3v//9Xrb9Y/HgwQOZTqfdzc1+xI3uVxCRTKdTARDG43GttcZqtZK6rrXW2hGR895nZ2dntizLbDab0e3bt0kpxVprq7W2nRNWe9C+0fsa8Mq6p7ve57Iftm2DhFf9I9gnDWLuDv39orOI2rS+6tbZVjmxS/vVZfStrrYFone3E1fHprixrQokbaNE4mYT0YwtRrSCPDNgTfOg9yDnmiXLgdEIMQT4GKGjNGHpsXPETyQSifek318GwROjZAXPCp65FT8YUAqkFBRRI3wAoBjAxiCOxvAHh/D5AJxnIOeaDKNB3lhdZRlgHcQYRKMRtW6u60YECUYjKt3YXREhEFrxo1nWGR/Aq4Bz3PDBicRrbE5g2yaAJHaLdruQiLCIaAC2qwAJITgRMUVR6DzP2VpL4/F4JzZiEkD2n25Hok0R4OHDh3j69On69ueff44//OEPP9jxvvnmm/V933///XvvmP/wD//wvk/56JyentK//du/XXUzrow///nPOD4+lv/4j/8AAJyengoA3Lt3TwDgH//xHwUAnj9/LgDw9OlTAZrKiPYH5dr3QbpA9KqqgrUWRCREpLXWcwAuhJBVVWUXi0XeBTlZa3MAA++9zbJMWWtZa325984NIYSAuq5RVRW89wghbB0k3BwYvG4CyC61/WOx+Z5+ysHdbdkd/XZ0nd+iKLBYLFDX9Xq9rgpkn8WCfph2/77+ZeLq2bZNNmep7du+l0gkPi7N4F4zw7qzxIIBYCzIOiiXgbMSVFeAD0BdQ6oSojSE6jSrJpFI/Cj6tlc1MSpWqEjBK90IIEoBSgNagbSGVgoQgdYaLBFwDuHgAOHgADIaIw4GTc5HJ4LkWVvpYZpFK0StEZRG1AqBGVFrRGYE5kbs4Fb8QBt23rW1Z3e1JvV3Ey39an8R+UEQemK3EBFqFxVj1F0ViIi4EIJFY4mlvPe8WCxoPB5fdZMBJAFknyERwaNHj+j+/fv09OlT+vrrr+nBgwd0fHxMp6entFgsMJlMCACGwyH993//9/rIcffuXdy9exfn5+ektV7ff3x8/Najy3K5fG0d59w7NXjzeR+Tg4MDrFarn/XIeHBw8HP+uTXn5+fr63meCwDcv39fXr58ieFwuO5XDIdDGY/HUhSFzOdzWa1WcnJyIqvVStr15dGjR/L48WN5+PBhBJpKiZ/9Df18dIHoAYAcHx9LnueF995qrefeexdjNFVVZbPZzIlIzszjqqqGi8XC3Lp1y00mE6uU4pv+I+y9R1mWePnyJZbLJaqqem0Q+scIID/VzP3LZm+/bd134afYD961DT92wPVd2rw50Puhf2fba2zLvOgLAl1nV2uNEAKKosByuYT3fut72Kym2PXv6LbPp1/9kSoLdoe+ALKtDD8JIInEDUcEQOuzD2qtZtrKEGMAo0HWNv75pQPZCmQNyFiQUmkAMJFI/GgimmqLmhgVKZSsUHEbQM4apBWgNWAMlHNNThERvOQgpiaT6OAQMpmARmNInoPyHOIsKMsgzgLWQLRpKjy4yTnyTBDV3W7sroQYEdIIIGgOjbIOZt8ifiQSW9gMPt/1c7obTheCrtsxNRtjtCJiY4xGKcV1XbMxhv74xz/Sr3/966tubxJA9hSaTqf05MkT+vzzz+n58+cMgP/pn/6JQgislKJf/OIXNJvNaDgckrWWVqsVHR0dUVEUBACr1Yq+//57AMB4PF7ff1lATV8kcc79YJ3BYPDWRvdf42NRVdVrr/ku7fhYiMh7vx+l1I/6DEIIrwkb3XVrrQBAWZZydHQkAOC9l8PDQwGA+XwuSqlIRNEYI3/961+jtTbmeR4BSFmW8eXLl72JGetB6OvaR5HpdCoiIo8ePYqTyYSHw+GKmXVZliaEYJRSeVEUeVVVw/l8Pjk9PR3eunXLAYC1VmVZpm/6D3EIAYvFAs+ePcPp6SkWi8Vrj7/vrPz3ESnel3e153qXdT5GBcvbPo/LHr9s0P/H8Lb3t21w/l3e57btuG1w+E0D/SICpdQ67NwYs36tsix/IID0BY99GoR+0+d5048vu8i26qSOfdrvEonEx0fQm8wBgbBqqkHQhAvDaJAxgNZQ1oKsBWkNUgpEaWZrIpH48Uhb+VG0wkfFGjUriDIQpSDt8Ue1OR2wFqIbuypYA3YONBwBwyGQ5+A8b6yveiHn0ehGUFEKNRECMzyksbsCWvGDEEUA6tldQRoVhHqB7InEJfQnRV5me5zYHboMkHbRImJa4cOGEGyboauUUmSModFoRI8ePSJcsfNMEkD2B5pOp/T73/+efve73/HR0REtFgsuikIxs/r00091CIFjjMzMqqoqHo1GHGNk7z0rpRgAteHPpJSi2Wy2vg4A3ntiZgKALqimw3u/vr058G+MQVVV2Pa8js37jTFvXH/butteU+vXd+GuHZc952MRQqB3PRB379EYgxDCa/e9DaWUAEBd14gxSndfXdfd60iMUdr11te11jHGKFmWRWaOdV0HAGE0GoXVahXquvZa6/DP//zP/uXLl+HLL7/0d+7ciffv349PnjyR1i6q679cO1qBR/7zP//Ta61LZtYiYrz3pqqqvK7rgfd+eH5+PqmqagJg8Ld/+7c6hPBu5U7XhBDCutqjy2FgZiyXS5ydneH8/Bzn5+eYz+c/qADZRRHkXV/3XcWGd329bRkV7/O33+V578Lbgpzf53Xedf1tllqXVTz0n6OUWgsgzAylFGKMl36W2yqQ9pWf8ruQeD/6+/qbLNsSicTN5dWgTetv31q/CDOguBE7tAJrDTCDlAIr3VSKpMNIIpH4WBCBtAbrxq5KjF2Lrpw5kO3yiBpxQ5xFzDJQloHyvBE7XCN6iHMQZyDWwqsmT8QrRqAmaD0ACJAm40MErZXE6yHnicR7cJkd8ub1xG5AjZc8D4dDe3h4mIlIrpTKmDkDYOu6NlprBUCVZcmdffVVkwSQ3YcA4OHDh/z111/zv/7rv/LR0RE/f/5cnZycqNVqpa21pqoqIyJaKaVExLSXipmV916FEFTr0cbee44xkohw67FHMUZiZvLeM/C6uBBjJCJCjHF91OmEknZddGrA5nrd85VS2LgPrfjy2nrbPgDvPTaf37bh0ud04cwfk82/1YkZl7Vh83nee/Q/07f9PWaW7n104oeISF3X0ntcmFmaVaIQURSRSESxvT8wcwgh1EopH2P0eZ7X3vs6z/NquVzWeZ5X3vv62bNn4fz8PDx48CCcnJzEhw8fypMnT15N4riGHB0dRQB+MBiUz549WxGRVUrNiqIYlmU5KstyZoyZ13W9DCEMAYRWPLkRv8DeeyyXS8xmMxRFsQ6i7jIZ5vM5yrJcZzN0bF5/kwBx2WM/96zqNw3qb2vj+3TC3kU8uaxS5WN+Du/6Gfc/i225B5vr/JgqkW0iSP/vd4JbjHFtg7Wt47RZAbIvneNtVTDbPofEbtFto/6++FN8VxOJxB5C6/8gBERqRJBIr4QR6gKJqT12pON8IpH4AAgCJQLdihDCDLEGsBk4y8DONVUezkG1YgfnOShzQLuIdY3gYc1aGAlaNyKK1q3w0VpdAQjUWm+B2vyRlO+R+HA2z3tS9cduw8xkrVWTycR57wfOuWFVVXlVVc57b733BoBmZrbWknOOvvjiC0yn0yttdxJAdpt11ceDBw8UAFZK6ZcvX6rRaKQXi4VhZrtYLBwzWyIyIQTLzBZt9F4IQTOzstaqGKNqRQ+OMSoA3IkfIsIhBGJmagUP6gbpRYS6ioVO6GgHQvtHo/Xj3cBA9/wuvKh/X/e6/cvN630uEzQuExJ+igPl5t/q/sbm/ZvvoX/be7/1OZvrElEnbICIpP28u/ukD4AYQogxxqiUiswcvPeRiCIR+RCCZ+YyhFBprasQQqWUKsqyLCFurlAAACAASURBVJ1zKwAlERUhBP/VV195a229Wq3C7373uwggPnnyBLimAsjTp0/l/v37wRhTlWVZEtGqrutFjHEmIjMimmmtF8aYpda6YuaPr6ztMGVZYjab4dtvv8VisUBZluvB6C4EHQA2K7HeVwD5OTo2P7byov/cbQLIxxr0fFerrvcZIO+3+11FijeJH5v3XSYavctn2V1/k4jSD7+7bNbIPtpfbbb1ss8ksXts+96n7ZVIJAD0Zj4LBIQQBRrt4CA1S7deOmokEomPAQHQEkERUKKgmUDWIAxyxHwAnedgl4HzV5UelLcVH84CziI6h6AUxJq18BGYGtsragLNAwQibeC6oAk5F2mObdvEj0TiPekmwG2KHkkA2U201uSc08fHx3mWZbJcLovz8/PBy5cvs8ViYb33pq5rpbXmuq754uKCnjx5cuUbMwkgu8drVlfffPON+s1vfqOcc8p7rwFY770JIZjVauWMMY6IMhFxdV07Zu4Hz1hm1mi2cyeAqL4AQkQkIkwtMcbuvm7npLZyhLpqkb7wccn1rYJG93xmhjGGB4MBZ1nGxhhuB7Be+0K8S5nUZYLJx2aj+uXSNmy+383nbluvv25fAOmLHv3b7XXx3seiKEJRFN57HwCEuq4jMwciCp0Awsy1974kopKISmYuiaggoqIsy6UxZrVarVbW2jLP8+ovf/lLba2tj46O6s8++yw8fPgwnJycxN/+9rfNOVyzma9FP+eLL76QR48exd/85jc+y7JqtVoVMcYVgCUzz5l5RkSzGON8tVot5vP5wFrrjDHaGMPMzBtC4LUixoiyLLFYLHB+fo6yLNfVWDHGtaDXeXR29Gfld7cv430G1n8qLhNh3kWUeFcRYhvbBIbNx973c3ibyLTtvb5JHNncFtteZ1vJ8mW8TQDpP3+z2qT9DXlrm3eZzcoX4JXlV57nYGZMJhPkeQ6t9d69v+uAiMB7j7quUZYlLi4usFgs4L1fV34mEolEn77nfTNTCQChGSBslygCgoBiBEkSvBOJxIdDbWWZUhrROcggh86HoOEQMhhCDQagTgDJcyDPQHkGOIfoLMS5JtxcawTFiFqjJkZUjMiMgKaCLbQiRxQBmBAltsc6uh6DAokrpX9O1E187s7/QghYrVaYz+cwxsAYA631VoeYxM8HEVE7jmu01o6Zs6qqstlsZkMINsaomVmJiFJKUZ7n9O///u9X3ewkgOwY1FldPXjwQHnv9Z07dwwRddUcDoALIWTz+dwRUbZYLHIAuYhkAJyIWBGxAGx73RCRFhFFRArAWvzoL53o0Q7mdgIIdcJE91gnYACvBus7YQPtEzbFjM3BfmstWWv1aDQyx8fHJssy3Q8H3yYi7AJvE1s2H98m6myu3398czC0Ezu6pbsPaCyxVquVPzs7q8qyrOq6rn0zGh2VUp0AEojIA/Ba66IVPkoApdZ6xcyrGOOyqqql1nrhvV9lWVYAKNvqkOLTTz+tnXO1c84/ffo0PHv2LE6n0/jFF1+s27LPEJFMp9OY5zlevHhR13VdxRhXIrJk5rnWeiYi50VRjE9PTwdaa1fXtTk4OMhGo5Fzzr0mCF43uoHAsixRliWWy+W62qO1oAMAKKVeO4nvBqrfNkjdDWpvEzzeNGD/vu/hbbzpOPM+4sA23tT2d62Ied8qize95jax4rKKj7dtg23PfdfttSlkvEls2vZ5bKtu2Ue6z8taC+ccBoMBbt26hdu3byPP89S5vwJEBFVV4eLiYp11dHZ2hrIsL93v9nkfTCQSH0bfF7UTPgSd8NFYOYYYQe11FmlmuYpAretFEolE4kfA3ASbuxw0GADjMfR4Ah6NIYNBU/GR5aA8hzgH5F3OR5MD4k0TiO6ZGwGEGZ6arI9IrcWVSGPlJ7HJ+ej67mivpwNY4gPZdm7aiSFlWeLly5dQSsF7j/F4jNFolM6RrphuAr21Fkop7b23WmsDwKIZuzYANBFxXdecZRl9+eWXV360SALI7kAPHz7k3/3ud7xYLLTW2mitLTNnMUYXY8y11pmIDLz3gxjjQEQGAHIAeQghExEXQrBodjorIgbAWvwIIbwmfHSVH+31tfjRW7Bx2Qkhr7W7N/DVfQ+w8dxNeDwe2/F4PLh9+3Z+cHBgtNbrEciemPIBH+fPz/tWo1wmfrSPvSYwbIoNIhIvLi6qGGPx/fffL7z3xWq18swcWpum2IkgALxSqmTmiogqZi6ZeaWUWjHzkoiWMca51nopIgsAK6XU0lq7ODg46ASR6quvvqr//u//3n/++ed48uSJSJM1svejPtPpVB4+fCifffZZ9N57EalEpFBKLQHMYoznFxcXw7/85S/u4uJCX1xcqF/84hcTrbWy1l77X94ugLq77O7bnLm4WbHwLt/fywbNN1/3Q44F71LZ8T7P/THrfKiAcZn4cNlrbz7+tkqN7jPe9rl3z7ls+26+3rsKEv3nd3/jXQSzd7lv19n87JRScM7h5OQEd+/exfHxMQ4PDzEcDlPn/groZpq9ePECX3/9Nc7OztYZSB2XCXeJROLmsXnCFAVQRGhjgQERSIyQGBFDAGIASWz7UVfR4kQicV2ISiFmOfzkEGE8RhxNgNEIPBhA8kErfGRAnkGyJusjWgMxTVB60ApBcSOAML2yvCIgAIigdWVbkzjS0EkgSfxIfGz655NdHmkIYe1Kce/ePRhj4Jzbu/HC60o3eb51HNIxRg1Aee+Vc46992ytpfF43I0nX1nvJwkgVw+hsb3i4+NjdXFxob33djweW+993oocg7quh8w81FqPh8PhRGs9ZuYhgCyEkMcYu1IjG2M0ImJERIuIEpEu7+O1pavo6NqAVuDYZnXVr1bYMuN9qyVW97zNN5xlGR8eHtrJZDKcTCaD8XhsjDE/EEDa1/uQz3bneZNo8qYDQwghiki1WCxWh4eHWQihdM7VzNyJErG9HogoMHOllKqZuVZKVURUaq2LTgQRkXld17MY40UIYR5CmHnvLREt67peVVVV5Hle/O///m99eHhYP3jwILTtvw4iiDx+/Dg+efIk/N///Z+31tbUZKKsjDHzEMJFURSDqqpcURSWmbNbt27ZEELeVltdK0IICCHAe4/VaoWiKBBC2Drzedss6Pedkf8u617lIOPHOAZd9hrvWx3yruu9SRR5k7hwmQi17b4PrYy5rH2dsLatGmXzNT+0Ougq2CYkiQiMMZhMJrh16xZu3bqFwWCAdkbNVTb3xuK9x3w+x+npKc7PzxFCgDEGSql1xdu+7XuJROKng4C1oNFdJxHEEBrhI0aEuoaqKshqBSkKoCqBGJBUkETiBkO0ttCLIKDrW/Tnk/bva+erUmt9JYMB4miCcHCIOJ4Akwl4MADyHJLnkCwDXCN+RKMRrEU0BlHrVvxQjdixFj9ay6tWwhU0t7tKj+Yy9X8SH5/LxhSqqkJVVet8kMPDQ9R1nfriO0Y7XqxCCDqEoL33WimlqqpSAHi1WvGdO3eufIMlAeRqoYcPH/LR0REDUEoprZSyMcasruusqqqRUmoMYBRCGAOYOOcOj46Ojkej0aExZhRjzEIITkRMu7OZVnVTIqL6YeftYDuLCAOvsj3Qm7zUHmjWl/22bg7Wb1nnnQQQay0fHR2ZyWQyGAwGeZZlr1WAJN5OjDGGEOrJZGJv3bpllFJlWZahE0D6IggaWyzPzJ6ZfXu9UkpVWusSwCqEMJvNZmeLxeJlVVVnAPKyLK333llrTYxRhxC4/Tvsva//67/+i/I8DyIS9l0EodYKC81klxpApZRaEdE8hHDeih/Oe+8mk8mwrutRjDFct9m/3UyLzu7q4uICy+US3vsfVBJ0l5szod/1M9lWPbKvvE/Fw7s8702fx/t8vpcJHpcJFJcJDN123iZ69AWL9/0+9J+z2YndDMHb3Oc+tDLoqtmsytFaI8syTCYTTCYTOOeuuIU3F2n9houiwHw+x2KxWG+nrvptc99NJBIJSHtsj7ERQUIAYkTwHlTXoKoClwVouYAqVuCyBLxvSkYSicSNpBE+AE+EQIxI/EroWC9t1iITmBXADFYKpBTiYIg4mSAeHELGE2A8brM+8sbmKssg1iI62wggulk6y6vAjNjZXVEbcg5pRA+0OUaxJ3rscd87sR9sCiHdxExqLYM7MSSxc5CIcAhBtxPxNQBV17UaDodsjKE///nPdP/+fZINt5ufkySAXCFt2Ln6m7/5Gw3Anp+fG+dcBmAwn8+HxphJWZaHAA5E5EBrfZRl2cnJycndk5OTk8FgMGZm2wkdMUZuhY9O8OBO4OiEiK6yo397o1k/sJ/qr/OmioX1C1zy3A6lFFlr1Wg0MlmWKWZOv6TvCRGRtVYdHR05Ywx/8skneQghto91AgioCVGPRNSJIaKUCgBCe5+PMZZFUVw8e/bsRVVVz5fL5ffe+9MYY26MOReRTCk1WywWhohW5+fnRQihqOu6+u677+ovv/wS10EE+f3vfy8PHjyIaDJTSmZeArhgZofGSs4ZY3JjzKHWumyra/b6PW/SzbI4Pz/HixcvcHZ2hvl8jtVqtQ7/3RwU7+5731kY+zCAeFXtuuyzfN/2XLb+ZqfxbYLLm/7uZQLGj2lfP/Suf982e659ZNtntOvfgZtKt526jKL+0j2etlkikehDRCARoPuNjREIARICoq8RywI0n0GfnUKdnUEvF+CqAsVwtQ1PJBJXhqARP0rWKLnJ4gAzhAmgRuSAYiitQUqBtQFbCzYGbA2QD4HRqBE+hkPQaNTaXfUqP7RGsAa1YnilUBMhMiGAEJjWlR7d2UEEGuu+9v4keiR+Dvq2yN3tbmHm12y59/Vc8LrSTazvLLC6SflEpJiZQwhcliUPh0N68uQJPXz4MFlg3TCoFT/0L3/5SwPAAciIKCuKYiAiIyIaV1V1qLU+NsYcZll2NB6Pjw8PD+9MJpO7BwcHt1sBxGCjmmND3NgqXlwmZLQHkw86orxNAGkPYmSMYa01pwPY+9POGObBYGCMMSqE0Ouj/CAvZB2k3j1ORBGAEJGEEGqt9Xi5XNrlcmm8966qKue9tyEE5713zOyIyAJYOOcW5+fnmohWd+/eJQD48ssvMZ1O43Q6Xbdj33jw4IHcu3cvfPPNN77NSym01gulVNZWZg2YeUREM+/9sizLYrVa5VmWgZkVM9NmBdS+0c2yWK1W6+Dfzvu+P9jXDVT/2OqPm8jHEi92gcva9rHavK0S5bqwTUBM7CZ98QPYD9E2kUj8/IgICI34IV3/KASIfyV+oKpAZYVQloirFVAWkKpKFliJxE2kq65AYztVs0KlNEqlUCsFsAKUAmkNKA3SGsoasDFQ1oKda5cMPBiABgNIa3uFwaDJ+sgconMIxsJrhWA0AjNqAjz6GR+AUHMY2jyJl2R3lfiZ2az87+7rxI89H2q51vQEENVVf3SLMYarquLj42M6OTm50o2YBJCfH3r48CHfu3eP0Xz+Tmudt3keQxEZi8ikqqoDETkiolvW2qPRaHTr6Ojo+Pj4+GQ8Hp8MBoOjwWAwZOa0DW8mpJQipRRb+2ExFG3wtxuNRlwUhQ4huPl87ubzuS2KIheR3BiTEZHTWmcxRgvAAOCiKAAAeZ7j3r17QUQC8Ob8kl1lOp3K48eP42KxCERUW2sLrbVaLBaWiAwzD5VS4xDCbLlczs/Pz+dE5EIIGAwGlojUdRFAqqpaW79UVfVaAHoSPa4fu7oNd7VdH8JllT2bNmOJq6c/42yzHL97vLtM2y2RuLm0wzUQiU3VR1cFEgNCVYGqGrGuQb5GXdVg70HeAzGCRVKGcCJxwxCgqb4gRq0YFWuUSqM2Bl5pQClAa8BosLFgawFrQa4RNShziFkOynOEPAdlGZBloDxDcA7IMgRjEK2B1xpBqUYE6YWbewhCV+XRXkLwuuCx36e1iT2lb3XMzK/ZIu+7BfJ1pZtELyLcRjB0WSCKmZWIqCzL2FpLn332GdDGpV1FW9Pg+c8LPX78mJ8+faoWi4VyzjlmHgAY13V9ICKTGONRXdeHMcbDGOOR1vq2Mebo9u3bx3/zN39zdHJycjgajUbGGAcg5WYkPhhmJmutPTg4mGitOcsy9/z582yxWGRlWY6892NjzMQY8zKEcC4iZ8ycGWOU1hpKKaxWK/zLv/xL/f/+3//Dr3/963CVvn4fwtOnT+X+/fuhKIpaKUVFUbAxxoQQDDOPROR8Npud/fWvfz1dLBaDW7duqTt37ggz02AwYObr8ZXcNusiDfAlEj+efkn3tu9SGkTfPfonWn3RYzO/JW23RCKxtgKV2FR++IBY1aC6bio9ihKx9ggE1NogWAcXIuABEwNUOo4kEjeG2IofhWoqPyqtUSuDaEwjfGgNMgbkLJR1UJkDWwedOagsA7WiBw+GkDwDnEO0dp310eV8BK0RFCMqagQPdFUfje0ViNZVa2hvJxJXDRG9ZtfciSDdY0kA2U3aChCWNggdbfWHUoq11myt5dlsxvhAt6EPJQkgPxPT6ZQB8GKx0CcnJ5qIDIBBURQTAEda6+PW7uokxngsIkdFURwOBoOjw8PDw1u3bh3dunVrcnh4OHTOGaWU3vfZ5ondgIjYGGOGw+FQa22Y2ZVl6c7Pz533fhRjnDjnDpVSEwAvQwgDZnYhBA4hQClFBwcHtFqteDab8dOnT+tnz57F1hJrnxKqZDqd4vHjx+H27dv04sULiAi16rVRSl2EEAar1erlt99+O7q4uMirqtLGGH14eNhVxlwr+lY9/YHANOCXSPx4tlkp9bNO0vfr6unPPNsUQkQE10XsTiQSHwHq/GMEEmJrf+URu+qPsoRUJUJdoQ4RSimI0hClYEKAxj51lROJxDvTWl01C62H/TwxKlYotEFtbCOKGg3Rpqn0MBrcCR9ZBp1lYOeg8hyqrfZo7K5yiMsQbRNwHk3zOnUbbh5YITK1AeeMAFmHnMfW3iplfCR2kc1hzq4fHmNEWZZYLpfI8xzWWiil1k4Viauhi2MgotdssERExxi1iCjvPX/66afriIZ2/Z/9pDcJID8D0+mUP//8c/7Tn/6kY4xmNBrZ5XKZxRjHAA5ijMfOuZM8z0/G4/E9rfUtETkuy3KcZdlkMplMDg8Px+PxeDgYDLIUGp74mFCDttZqpZQJIZjJZKIPDg40M+cxxpFzbklEwxhjvlwuTQiB0diGhhgj6rrGcDgkrTV99dVXCCF4AJhOp9g3EeThw4fxyy+/DLdv38aLFy+6fA9jrZ1XVTVfrVYX3vuzxWIxtNYOTk5ORt57jz3NPnkbbwptTgO1icS786Zw+76dUmI36Isgl+XSpO2VSCSayo82/6O1wJLgAe8hVYVQVYhVBdSd7RXAxDCsEKjx308kEtePuF4IkRnS9hm8UqhYozIWtbXw2gBGg5wDWQuyFuwyUNaIHpRl4CwD5zmQZ6Asg+Q5Yp4hWItoTBN0rhUqZnjm1u6KIOu8kVb8kFeCTMr4SOwq/cliXQVIZ9U9n8/RZrBiNBphMBis++uJq6MVqBiNSxGLiAKgtNZKa83GGJ7P510FSLLAusYQgLX4UVVVvlqtcgAjIjoAcNt7f1trfffg4OCTX/ziF//fcDi8bYw58t47IsqzLHNHR0eZc06nk+3ETwkRUZZl6vDwMCMi1HXtRGRkjKmqqhosFov8+++/V7PZjMqyFKUUyrJUWmsVY1TeezUej6ksS/rNb36D+XwuV6Xu/liISKbTafz8889x+/ZtrFaryntfiMjKe79QSs1DCHOt9VwptdBaF8wccI0EkDcdZ5LlSyLx/lwmfHSX6Tu1W/QFqW3l9tvC7FP/LJG4oXQ5Hp0QUtcQ74HW/krqJgOkuw3vEUKNGHxz/EiH/0TiWiJ4Ve3hmdciSFAaXil46xCNWYsecE3FxzrkPM+bbI9BDmQ5YubavA8Hca4RP5xDVM3rB9WIH56osboiQuzyPYjWmR8grLM/Ut8lsYts7pudCLJcLvHtt99iNpvh7OwMn3zyCU5OTjAej5MAcsV0VSAxRo4xqi4LBIASEcXMpJSiP/3pT/SnP/2Jfvvb315JO5MA8tNC0+mUjo+P1bNnz4xSymVZlocQxjHGAyI6NsacMPPd0Wj0ycHBwb2Tk5O/nUwmt/M8n7Q7jWZm5ZzT1lpOP1KJnxIiIq21Go/H1lqrYowZEQVmDqvVyhljTFEU4r0nEYnGGGFmqqqKiAhKKVqtVsjzHFVVCQB58uQJRCTukwgynU6jiMiTJ08EQK21rmKMhTFmSUQLADOl1EwpNY8xruq6ruq69kSklVLU/gDv9Zf1XcLGkhiSSLydy04w+wPoSQTZPfrHvm2l+P3radslEjeUTgxtKzsQGwsseA/piR6xqiBVBfIewdeQEBpPcxFIUkASiWtJpCbro2INrxvRIzIjKoWoNaJpcjvgmoBzyvO18NFVfHQiiOQZxFpQ3lpeWYtgNKI2iKoNOGeCJ8ATratPpMtT6FV7dKHnaVwpsev0++Gd68h8PsfFxQVWqxWyLMNkMsFoNLriliY2BRAiWosfIqK6HBCtdcoAua5Mp1O6d++euri40MPh0JZlmYcQxiJyKCK3rLUnxph7zrl7t2/f/uTk5OTe4eHh3clkcpjn+QhodiQgBf4kfh6ICFprVkqxc870w8yVUjrGqIqiABEpay1CCExEKoSgRATeezLGSIxR7ty5E8fjcfzqq68ArC1Q94b2fYfHjx/7ly9fVnVdFyKyAjAPIcwBzOq6ni0Wi8Xp6enKez8YjUY8GAy0tZb31apuM+Q3DewlEh+fy6zlErtBX/ztLLAuC0BPfbNE4obSff9jbPwcRBoLrBAgdQ2qauD/Z+9eliQ5jvUA/+4Rkbe69XUADHlAUXZ0sYG04koLGbngRg8w5xHOa6DnGbTSeQRiqwfA2WjHJWAmk4ymCwQSBDEzfauqzIhw1yIza2qaPYPBjVXd7R8tUTXdg0H2JDMqMjzcfQh89FkhEUgRlDMkpU25rLs1OzbGvCsF9VkZ3qPzAdF5iOO+0Xno+31gyPag+lXAYzxoKHmlVQUt+9+rQ8mrHPom52NmiWAMuABJdVP6SlWhN0t5Et3tXXrm3tveXLS9YSzGiMvLS6gqRASPHj1CjPG1pulmd4bgxyYDZAyCjI3QxyyQXWV/ABYA+cmoKj179oyvr699Sqnouq5yzjVd181yzodEdDKZTN47Ojr62enp6c+Oj48fzefzk6ZppiGEgoj6LeT2YG3+tjYBt61XAoCiKIrJZDJVVW2ahi8vL3F+fk5t29JqtQIzpxCCpJTy1dWVxhilrms5PT3VTz/9dOwZcuecnp7K119/nVU1OufWqrqKMV6LyNXl5eXlF198cXFxcXF5fHxcPnr0iD744IPKORfuehrm23Y/G2O+u+3F8pulkyyLYP/cbIJ+03YJMxsjjXm4NsWsJYNVQCJ9v4/YQWMHyhk0NEbHJvihm8bpxph7igigPuChvm9yTqEPfqj3fTmrsgBVNbipwE0DqipQ0wBV3+RcyhKoKkgRoEWfMZIdI7uxrBa9am4+xFMFr7I8ANtkY+6ebysvaxn0+2nYvD8ejD4DhEWEvfe8Wq348PCQfv/739OvfvWrnZyjBUB+GvTJJ5/w0dGRAxBSSiWAWlUnqrrw3h8x82nTNO8fHR198P777z9eLBYnk8lkUZZl6Zyz62L2jnPOV1XVOOd8URTOew/padu2AiCmlARAds7p5eVlds7li4sL/fu//3s5OzvjO9YQHQDw9ddfa9u2+eDgIK5Wq05E1kS0TCldX1xcXL18+fIqhHD53nvv1aoaFotFaJrGhxB2feo/yPYO6O3dzsaY7+5ti+TjLiazP97UA2Q7E8TGQ2MesHEswPCkPwY0cgal1B8xQruh70eMfWZIzmARkEqfMdL/YTv8QYwxPxkiwDHgXN/YvCihvn+PogCGnh5j9gdNGnDVZ3702R81tCz6fh8hQIuA7Fzf8wMYen302R6iCoG+iqnaPMXcE9tz7+2NSTezs83OkfeenHMuhOBzzg6A40GMkYuioLFKyrNnz3bSCP1ub1HeT3R2dkaff/65W61WxeXlZQ1gklKaL5fLw6qqjmez2aOTk5MPjo+PPzg+Pn5vsViczGazRdM0E+99MaQKGbNXiMh574u6rpumaeZN0xzPZrNHs9nsvel0+n4I4TTnfNx13WHbtouu62aXl5fNfD4vv/jii/DrX/+az87OGHesN8bnn3+u//bf/lsRkey975h5TURrEVleX18vnz9/fv2nP/3p+uuvv15dXFx0Mcasd3jGub2T4uarMebHdfPesntt98aHqjGL77ZgiD10GfPQ0WtbHBkKpwonCicCHgIgHCMoRlBK4JxBImBVUF+bZvNnGGPuISaQD6ChublvGvjJBG46HLMp3GwKns7A8xloOgVmM+h0Ap1MIHWNXFVIZYFcBCTvEZ1DZEZkRiIgEyFpnwEylrwS2xVv7om3/f/Y5uF7hZxzXFVVmM1m5cHBQTGbzYrpdOqcc05EOOfMbdvy8+fPqa5r+vjjj3dyopZp8OOip0+f8gcffMB//OMfC2au67qeLZfLAyI6TCmdFEXxwenp6c9OTk5+cXR09P7h4eF70+l0VpZlZZkfZp/RAAAXRVFOJpMZAPXeu6IowvPnz6VtW7darRwzh6IoSERovV5TCEHLspQnT57k3/3ud/kf/uEfxnnanXB1daXz+TxfXl6m5XLZDQGQVYxx1XXdSkTWMcYu55y0t+tT/sHe9DPch5/NmF14U7DDAo37Z3ygcs5tdpuNbmbz2MOXMQ9P3/NjCIBof5AoKGdwTH3z87aFdh3ckP0hOYNUQdIHS2wXojH3GxGDvIerKuikD2qMfT9QFtCmhlZVn+lRlUA9lLwqS8iQ8SE+IHuHzAwh6vt8QCGgV0EPDHNIIuvvSfLpxwAAIABJREFUYe6Fmz1A3nRYGdr9wMxUlqU/ODioiGiyWq0m6/W6Wq/XoW1b55xj59ymB0jOeWfnagvuPx5++vQp/fa3v+XDw0N/fX1dtG3bqOp8DH6klE699+9Np9MPHj169LODg4PTyWRyWJZl4ZyzrA9zZzCzL4qiISLvvXfM7K6vr7sQAkQEREQiIjFGHTIikqqmuq7jarXC7373O9ylIMiLFy/Uey8hhKSqMaXUiUirqmtVbYmoc85FZs7MLGPj+LtmO710+7CJhTE/ntvKJ1nwY//cHA9v7jT7tvrExph7ShU0ZIA4ADxkfrAqKAsovmp+LmMT9JTAqtAhC4SGAIiNHsbccdtzgM176m/uEMBliTBpwLMpZDIFVRW0KPq+Hk0NGQIfuSwgZdmXu3IOEjzE+z7w4dwQ/Bj6e4D6clfYepC2uYi5Z27bbHSz54fNwfcDM1NRFG6xWJRVVeW2bSfX19fV+fm5v7i44K7rmIiImTclsHbFAiA/Dj47O+NvvvnGXVxc+Jxz4b1vcs7T9Xp9oKqHKaXjnPNJzvnUOXdS1/Vh0zTzuq6b4f8EthHI3BlExN77wMwegIqIzmazNuesIoIYI3LOKeecAEQiit77NJ1OCQDuUhDk448/1k8//VSvrq7yV199lUQkElHHzC2AlojWzNw65zrvfWLmO13M3zmHsiwxmUwQYwQzI6UEEbFFWmO+JyIag8OvZXzcXES3e2x/3Nxltv1164tkzAM17jYdgiCsChYB5wy36f2R+t4fbQd0HZDS0ABdNlkjTocMErUgiDF3nRJDnYN6DzgHJQI7BuoJaL4Azebg2RyYTPreHmU5ZH5UfbZHVQJFGHp9eCTu/7zMjDxkfShT3+sDQ5kr9Bkfr2V/GHPP3Jx/jxuTxgwCa4K+H4gIQwksCiEURVEUzBxWq5VnZsfMnHPmMQBSFMXOBiwLgPxwNPQ18HVdhxhjsV6vqxjjLOe8EJHDGONxSuk4xniaUjpKKS2IqHHOWcNzcycNpbCccw4hhKosSzk8PIzee4QQ+OrqSq+vr7vVatV57zsR6bz3MaWEqqr0+PhYi6LQs7MzPTs72+tPLSLC7373O72+vpbcj9xpKHfVMvMY/Gidcx0zJyK60xkg3ns0TYPj42M453B5eYmrqyus1+vNJMMWa415d7elaN+Wsm3NtffHdtDj5uv43q6TMQ/MduNzxaaRucsClxJcTEDX9/0YMz/QddAY4USAIfODdOwbYsEPY+48oj74UdXIdQUtSsAHiHeQZgKZTIHFATCdgiYTUFVCyz4LRKsSOmR+5OCRQ1/uSobARyb0pa6IoDTsGByzQIYpiAU/zH30tuek8T2ATb8+s3M0XAvi/g2v12vnnGMiYtoy/guffPLJTgYuW3z/Yejp06f8zTffuOPjY39wcFBMp9NaRCY553nO+TDGeBRjPI4xnojIyXq9PmzbdppSKkTE7lhz5znnfFVVNREd13XtyrL0ANJqtVqllNbM3BJR65xrvfdSlmVeLpeyWCzkyZMngv75b+9XkiaTiSyXy7xarRKATQDEObd2zrUhhM45l+5q8APoJxNFUWA+n6MoCpRliRACUkqbwxjz/dzWO+JmRojZvdtS7rcfuqz0lTEP0+aeHwIYpABngcsZPiVQF0FdB+o6oO36LJAugmMC5QxIBqmAMZTO2uHPYoz5kRBBvUeua+SDwz7gUVZACEDTQOt6k/mhdQUdSmBpUUCKAlKEIfjRNzjPY7krABlAHjI95FXEA5tSAzZvNA/AbYGP8b31ANlPqkoASER4NPYAuby8pLqud3ZuFgD5gT766KOxBGzhnKtXq9WMmefMfBRjPBaRE+/9adM0p2VZHp+cnBzMZrPJUD7I5r7mzhvLYRGRA6CTySSHEC6J6CLnvATQqmrXdV0MIWhKKa/Xa/nDH/4gL168kDuQBaKff/65fvnll/r48WNp2zYxc6yqqr2+vh5LYK1yzqv1er16+fLlyjlXTadTLsuSh6ZPd+KTeUhf3AQ+cs5Yr9coigLWpsiYH26cqL+pFJbZDVVFSgld12G1WuH8/BzL5RI559eukz1kGfNAjbust0pgMQROMnhodE5t2x+rFdxqCVxfQ66voKtVnw2SIiglsGR4FQRVOKhlgRhzFxD3ZaichzoHONePCc5B6ho6P4AcHkGnM0hVgash2DEcMpS6kqLom5uHgOR93+DceyTHyM4hMyErkFX7kle6leUxzBcVtgnD3G83y8+OX9t+NftrDIAQEYsIq+qmBwgA+uKLL6wE1l10dnY29u7wTdMUAGpmnqaUDoZSV8cicjyZTI7m8/nR0dHR0fvvvz87Ojpq6rr2FgAx98FYDst777z3JTM3IjLLOS9yztciss45tymlVlWjiHTz+Tyen5+nv/u7v0uHh4d7nwVydnamT58+lX/37/5dXi6Xab1ex5RSVNWOmVtmXsUYV+fn58svv/xyGWOsDg4O+OjoqGiapq8VdkeMDX8BoCgKeO9fm3DYQq0x389tDbS37ye7t3ZHRNB1HV6+fImLiwu8fPkSl5eX6LoOAGwMNOaB24wBQB/8UAVnAacElyK4bcFdB1qvwasVeHkNXF2Crq+g6xbataCcQdJngnhVBCjYAiDG3A1D8EPqGlKUQFkCzgPeAXUDnc1BB4fQ6RRc10DVNzTXsoKUQ6bHkPWRfZ/pkcc+H8zITEg0BD4ACKFvc04AsDX3GMrwGXPfvcvGIwuG7KfhuoxBkM1r27YUY6SyLC0Achd99tln9NFHH/F8Pvdd1xUAGlWd55wPReRYRI4BHFdVdfzo0aPDDz/88ODRo0ezg4ODajKZBO+9BUDMvaKqnHMOOec6xjjPOa9EZK2qrXNuBWAdY1wxczufz2POmeu6prOzM9rzLBB89NFHWpalPH/+PANI3vvonOtEpCWi9XK5XP7pT3+6ury8vDg/Py9+9rOfcVEUHELgEMKuT/9HYTugjfnhbAF9/4gIlssl/vKXv+Crr77C+fk51us1cs4Q6YtNbAc/bBw05gEaM/hEQDI0P08JLka4rgO3a1C7hl8u4S4v4S7PwZeXoBghKfX9P0ReBVCgcLA+IMbcBUoMDQG5mSLP5pDJBFwUoFAAVQVqJuDZDNTUQ8ZH/3UtCkhZIHmPVAQk7jM9EnPf42Nocp7R9/aQIfMDwKsG58Y8MLf1Tvy292b/qCoREakqp5QohEDz+RwvXrzA06dPd3JOFgD5nlSVnj175k5PT/3Lly9L732dc57mnBfOuUNmPp5OpychhOOTk5PD09PTxaNHjybHx8dVXdeF956HFCBj7g0iYuecL8uymU6n85RSVxRFq6rx+vp6TURr7/0yxtgSUZzP53G1WsmTJ090GCD39VNMz87OMARppCiK3HVd8t53ANYAljHG64uLi6urq6tL7309n8+LGGMpInd6nL0tBXX8OmATD2Pe1W3lr7bZovruiAhijFgul5ssEBGBc25zzW57ELNrZsz9tr0Iw0R903OgD4LkDIoR1HbAeg2s16DValMCK6xXcO0alFJfQksV/YbuYfzYOowxe4IIygxlB2UGiEGuD35IVUMODiDzA+hsDikKUFmAqwpSVkD9KvihZYFcFsghIBWhL3PlHSL1GR+J+iwPAUGgr4Ifw2nY85V5yLbXGW4+O23Py60s1l4jAJsm6EMrENr1GvidXpjbFVWlTz/91H3wwQf+m2++KUWkSilNUkrznPNhzvm0aZpH8/n80eHh4enJycnRe++9Nz88PGym02kRQrC/d3MvOecohBDm8/kkpRSLotCu63KMMccY1wCWKaXrsizXzrlutVp1dV3LL37xC8Ww0WXHP8LbKAA5OjrKYxZIWZYtEa0AXMUYL1ar1STGOFksFpO2bWsRmeg9mcHaxMKYH+a2wMfbgovmb0dVN2WwVqsVVqsViGjT/2gsC2glsIx5WGgoN7MpfQWAtM/+oKHxua7X0OVyc2C9Arct3NAbhHPe7Q9hjHlnygzxHrmqIb4AhQD2HijLvtfHwRF0voBOZ0BdAUXR9/coArQo+/4eRUAOAXkIfOTgkJxDIkIkgjANDc7Hh99+bmHNzY153c2m5zfZnHw/qSqN2R9jI3QazGYzNE2zs3Ozhfjvjj755BOeTqcOQJjNZuX19XWzXq+nMcZ5SunQe38cQjg5PT09+fDDD08ODw8Xi8WibprGGp+be805x3Vdh6Ojo6YsS51Op/zixYv08uXLuFwul0R0GUK4aNt2CaAlorYoinx+fp4//fRTGdJA9vaT7OzsTP/Lf/kvUtd1Xq1WiYi6oihWKaUr59yl934mItfe+xUzd0SUmVm+/U/ef+MOjNt6FxhjbvemTA8R2Sy62720P24r8/emRox23Yy5/8bgB4/vx/JVQwBE2xa6XkNWq77Z+WoN17bQFPuSWbs9fWPMd6TsIEWJbjKDNhNoVcOXJaiuQHUNnUzB0xl00vR9QIoSeWhqnovQB0+8R3aMHHyf7cHcl7kiQoYia1/uSoe5xL7vADRmF27OvS17/m4YAh8AQCLyWg8QIqLr62s6Pz+nn//85zs5PwuAfEdnZ2f04sULXq/XXkRKVa1TShMA86qqDpj5qGma49PT0+PT09PDk5OT2WKxaIayV27XKT/G/JSIiL33mEwmxMzqnEPOuUspxZzzMud8DuCliFx1XbcSkXVVVVFE0qNHj/KzZ88Eez4H/OMf/6iTyUSm02m6urqK3vtVCOFaVa+HQMg1M6+ZORLRvQl+GGN+mNvKxo0L6XaP7YebafU396zcvHbGmPtt+55nACQ69ADJoJyhsYO0LdC2oHX/Kl0HTQId+n0YY/YQc99rgxlKDBABBOSyQq4byHwBnc6hkwlyVYKrvrE5mgbaNNCq6pucF0ODc+8QnYf4obG5225u/qrMlRL15a6A1zaVKdCfgzEGwJs3Jd1k8/H9NGSB8HjknJmZaTqdYjKZ7Oy8LADyHX322WcEwD169KhwzlUppUZVp977WV3XB7PZ7GixWBwfHx8fHR0dLRaLxWQ2m5Xee/u7NvceEZEbMDOYGV3XpZxzUtVl13XP1+v1XETOVfW6KIqy67rWex///Oc/x48//hhnZ2e7/jHeRj/77DP9D//hP0jbttl7H7337RAAuUopXeecl8y89t53zrkxu/nOsoVZY34ct91L1shvP9wW+LgZBLl5reyBy5j7j4a+H2PzcwbAOgRCcgZShnYdZN2C2hboOkiMkJygYmO6MftKiSDeQ32ftQHnASZo1UCaCbA4hExn0Om07/FRV6CqhFYVUJXQsoKMmR9h6O/BDuIYiQiZx+bmigyCUl/yCuh7ffQBF7LghzFvcLP33psqUdhGsv1zMwsk5zxmguD6+pqsBNYd8tvf/pZTSl5Vy+VyOVHVmYgsqqo6PDo6Ov67v/u7RycnJ+8tFouTyWQyq6qqICIre2UeHGbmsizD4eHhtKoqnc1m64uLi29evnw5Pz8/n4nIdc75uq7rFkA3m81a3IFekB999JF672WxWKRvvvkmOuda59ySma+H7I/rEMLKOdcx870pgWWM+XG8rRG62a3byl2NXx+J2JBuzIMjfUYHKQAVsCo0ZSBGaBehXQcaDo0JyEMGiDFmL6lzkKJCHMpcoaoA7/v3zQQ6nYKaCahpQHUFVBW0KiFF0Wd9lCWk8BDvkTwjsUNyjAgMgQ/0WR/EyEPAQ4aFWiLqy16p9lliFvww5jXbzc1VFcxsWdh3zNgHBEP5KwxvdnxaFgD5LlSV/vN//s/svQ9EVKnqJOc8V9UFER2UZXmwWCwOjo6OFrPZbFZVVRVCsLJX5kFiZnLO+aqqyDknzrlZjHF2eXk5VdUJgIaZ65zzajqdrsqy5E8//fRO3CvPnz/Xtm2laZoIoBWRdQhh2XXdkplXzNw65+5NCaxttvPZmO9nnLiPk/nt8lcWDNm97ety22HXyZgHbJz7SO6DICIgVSBnaM5ASkBMQ/Aj98GSu50AbMz9QkNHH+a+0XnZ9/PAdAZtptCmAYqi7/NRVqDpBKhqoK6hZQEMwY9Ng/MQIN5BvEMaS10xI6EPgPRlrrQPeowBj+E8ZJxLDFkgxphXbmZ73DYHt+enO4O2dV1HOWdqmga7WvezzIR3pKr07NkzKsvSEVGIMTaqOss5LwAcENEBMx+UZTmbTCaTIf5ROOfcPkS6jNkBds65oiiKqqqqoiiaEELDzBNVnYhIIyK1qpar1SqsVis3m832/l45OztTAHJycpJDCGkymbRVVa2GxucrAGtmbokoYijxutsz/vFYA3RjvrvtXUzAm0th2X21W+MOs9F28GPbm7JEjDH3E42LlONijGofABkOTRHICZoSIHnzen9mf8bcE8xQH6B1A0ym0OkMtDgEHRyADg5Bxyego2Pw8TH44AC0mIPmM+h8BplNkacTpKZGrErEskBXeHTeIXqHbmh2npn7ZucEZOrLYI0BkTEQYoEPY97utrKzNwMh9ty0v8aEDwwlsMZm6GVZYjKZ4Ouvv97ZAGgZIO9AVekf/uEf+Le//S0DCCJSdl036bpukXM+EpGjGONRjHExBEb8kO5jjBkQEYtIkVKqRaTJOU9EpI4xVgAKInKLxYKGmoF7/Yn25MkTBSDOuaSqUVXXAFYAlkS0JKKWmaNzLu/7z/IubLHPmB9mO3PqTc3Qze5t7zYbX28+eBljHo5xsWXYOz4cunmVMRNEFQSF5qHxuQIWATFmjxBBvYc2DWQ6h84X4OkMPJ312R/NBKgraF31Dc7rGlSWyEUBLQNS8EjOIQ1NzTcNzoFNU/MsMjQ5HxZox8PmDsb8IDfvIeuhuN+2yl+NPYIBAF3XkYjs9KHXAiDf4uzsjJ89e8b/8T/+R3dxceFDCFVKadK27Rx95sdxVVUn0+n0uCzLQ2ZuVDXgDvQyMOZvRVUp5+xSSkVKqc45N6radF3XEFHFzMX19bVr25afPHmy69P9Nvr555/rr3/9a/lf/+t/5aOjo+7Pf/6zTymtU0rrnPNaRNYxxna1WnVFUUQiSn1feKa7WhJve4HWFgKN+e7eVj7OdjPth5vj3G1fs2tkzMOxHfgAsCl9tTkw7EbNQ0aICqDbQRBjzE/iRlmpYfvC5p+k/XeJqM+88B5aN9DZAnp4BJ0vQNMZ3GToAdI00KrsAyB1jVyW0KHPR/RuaHLOiFBkAIkISWVT6mr4r0FVNre+DQHGfH+3zcNvsjn5fhsqIW0aoe/6fAArgfVWZ2dnjP7vyD9//jw450pVrYfSPTNVPQghHC4Wi6Ojo6OjxWIxL8uyds55K3tlzGsIAOecQ865FJE651yJSKWqBQBfFAV//fXX9OzZs9eeNffR2dmZ/vM//7NMJhNh5tw0TUdEnap2qtp1XddeX1+3z58/b1++fNleXl7GGGMWkTv9KW2lX4z5/m5mftxcTLdJ/H74tjHOxkFjHpbNIsz4fhiqNw2MRTav2wuvtvxpzE9HAQgImRiRGNH5147MDCWGMENCgNQNZDqDzBeQxQH0oC99hdkMtDnm0MkU0jTITYNcV8hVhVQWiCEgBo/oHJL3iBiCIMzIwHDopvax3f3G/Di2N4lZyeC7RURIVUlEOOfMRERN0+C9997b2TlZAOTN6MmTJ3R0dOTqug4nJydlWZYTVZ3FGBfL5XJBRIvJZHLw+PHjo1/+8pdHH3744cHx8XFdlqUFQIy5QVVZRHyMsYgxFkMgpBCRoKrOOUd1XdPHH3+861N9FwoAp6en8pe//EVUNTNzApCIKF5cXLRffPHF8r//9/9++T//5/+8+vLLL5dDEOTONkW3yYYx39/NZn7bpZXGr5nduZmBc1smyM33xpiH4bUFl5vZepup0evfh82ZjPlJKfoeG63zWIUC16HEsqqxqhq0ZYXoA7Jz0FBAJzPkoxPkk0fIR0fQxQKYzSDTKWTWH6mp0dUlurLA2ju0nrFmwgqKDkAHRVRBUkUSeRXoELEyV8b8BG7r93GzJK1tStpf43VhZowlsGKMO79YFgB5A1XFixcv+Pnz5y6EELquq0Rk0nXdLMa4SCnNRWRRluX8+Ph48f7778/fe++96XQ6rYqisMbnxtww1AJ0IhJSSmXOuVDVICIhxuivrq5cURT0ySef0F2YRH788cf69ddf62QykfPzc8k5ZwBJVdPFxUX805/+tP7DH/5w/b//9/++/uqrr9bX19cp53wnAyB34XoYc1dsaspvTeDfVh7L/G3dfOASkbc2sDfGPAT02rbuzfhNr8rtkPYlsGhTJgu2DdyYn4iiL22VmRF9QBdKrIsSbV2jqxrEskIuSkjdIM8XyIcnyMcn0KNj6GIBmU6hkwnytA9+jM3N2yKgKwLWzFgToSNCC0WniiiCDEVWhUAhqq+CHzaHM+YntZ0BYs9MdwMzY7sJOgCsVivrAbKPnj17Rt988w3//Oc/d6vVKoQQqhjjNMY4jzEuhgboMwCzpmmms9lsslgsKiJiuyGNed0Q/GARcUPGRyEiZc65SCkFIvI5Zy6Kgp4+fbrr030nRISzszP99a9/LS9evJCUUlbVBCAtl8supdSKyBLAarFYtG3b1jlnexQ2xty6q8ns3riTbFzcvBmoMsY8TIQbi5yqYCKI9l9nAJwzXErwOcOJgKwQjjF/IwRlhlYVJBTITJBYQVSAqoQsDiEnJ9DFAdA04KYGmhpa1X3D87IY+nx4RGYkx4jMyIwh4AFkVSgNDc+HwAdgwQ9j/ta2AyFWEms/Dc9Sf1XWPsZIRETffPPNzgZNywB5g88++4yOj49ptVq5GGNIKZXOuSbnPM05z1JK0xjjpOu6OqVUAHA0wI1+ecaYV43Qc85BVUPOuRCRQlUDABdC4BACffrpp3fl3tExC6QoCokx5pxzVtWUc04AoqpGVU1DYORePQlboNeY72Y7i+Bm+vb2q/nbu/l3f1spLGPMwzQGP/r+H6/3bVJVsCo4JxQpooodqtjB5wQeeoIYY358hP7eCzmjlIyKFMF7cNMAiwPI6SnyB4+R3n8Mee89yNEhZD6DzmfI0wlS0yA2FWLdZ33EskTn+4bnnWMkJkQiJCJEDD0+VJG3y18BFvww5ifypgCHzc33n6puLtJY/goAiqLYyflsswyQt/jyyy/5+PjYOecCM5dENAZApimlaUqp6bquyjl7EbFgkjFvsVUCyw9BwyAiQUR8ztkTEV9cXNB/+k//CRieN3d7xt+OiPTs7KzvwwdISimLSGbmlFJKRDQeQkTjfNkY88DczCjYLqtk9s92Jsj4aytXZszDM7Y/J0Lf7Hz8miqg4443BYsgpIQyRhRdCycCtl2pxrybrc/U7btm89XxXhp/HxGIGEyEQAAz4LwDVyXybAqZTIGiQC4CuKqhdQ2dNNCqBqoSWhbQsoKWJaToe4Uk5r6pOREiaR/woD7rY8zfVyLL/DDmJ3Zb772bWfOW9bH/xrJX4+tYAqtpGvSV43fDAiBv8NFHH9HV1RXFGJ1zzrdtWzJzLSJNSmkiIvWQ/VHGGL2IsKpa6w9jbjFEgWkogeVFxBORH98PgRGu65p+//vf0x/+8Icxi2rvP93Ozs70H//xHzWEoFVVCRFlEcnjK/pNQ3ey94cx5sezPVm/uaBu9sObrsltv7ZAiDEPx2tjgOqwMDuMF6JgBZwIvGR4C34Y851tdpNtwo4AQ18vq0EEZQf1HggeYAdihisroGmgizmwmAOzOVD35a1yUfZlsIoSWoQ++BEKSBE2wY/MjMyMRH1j9aSKDOozPVT7fiNQqOhrQRhjzE/ntk1I29+zOfj+ExECQNtZILtmAZC3YGZWVUb/91SsVqsmpdQMmR91jLGIMQYRcdtpPsaYv6aqmwCIqnpsZYCklFxZluy9p7quh811d2ZxSR8/fqzr9Vq6rhMAQkSbclgAMjNnZrYgiDEP2G2NtLfHOatju3vbD1vjA9f255BdH2Menlf3vW7KYSlelcbi/jf1fUCGkliwscKY70QARGJE6otqOFUEFTjoJgCi7CBF0Tcwr2qgqkDeQ6sKPJmAFwdwsxloCICgrqFFAQkBWgRk75GdgwSP7BjifB/8AJCZ+ubmKhDq3+vYyUelD3jcjedSY+6dm8EQKx+8/5iHsdw5pJTIe4+yLHd8VhYAeaMvv/ySDg4OEGMkZvaqGrz3ZYyxTinVKaUypRRSSi7nzCJC9mBszO2GDytmZnbOeedcUNVARB6Ac86xiLD3ngDgrjRCHz158kT/23/7byoiqqqbIAiATESZiET7FLF7MUjcoeCUMXvhbRkFlgmyX27uKhMRMLNdH2MeKnq1A13Rz3/6nTpbzdGNMT+IgJCJ0DFDAXjtM6tYFaA+5KhDsCPPFtD5HDqZgssSqCtQ04AmE/jJBDKZ9GWvqgo5BKj3yN4hDdkekQjiGAmA0JCqrwqFvsr6GEuXAhb4MGaPjKWEAVuT2HfMDBEh5xxyzntxoSwA8har1Yq89xxjZOecyzlvGjePO9ct+8OYd0Lee67rOszn81JVq5RSMQRD3Bj8cM5RURT06aef0m9+85tdn/M7+/zzzxUAnHMqIppzFlWVIevjXgU/RvbAb8y7eVP5JLN/bsvSuZl6f1sqvjHmgVEFEaBb9XlsbDfmR0IMZUKmfgFNeci+qGvIZAo5PITMF8B02meBNH2wA3UNqSpg0vT9PcoSEvoyV5FpKHM1lLoCkKAQBQQKoVeJW33Wh93LxuyaBTfuLhGhoQTW3gQ/AAuAvFXbtpRz5qqqWEQcAK+qfmh67nLObrywFgQx5s2IiMqydPP5vBSRejKZ1Ov1ulytViHn7HLOTES0XC7v7H20XC61LEsFoESkRKTSb0/QoQH6vZtM37efx5if2m2ZHzffm93ZXsC8mQlimTrGmNf6EWDYfdq/wx1oW2fM3iL05eO8CNQzKPQkx5ZHAAAgAElEQVQ9OqIPcEUBeNeXtJpMoYdH0OkMNJsilyWoroCqghYFtKogZQEp+ybo2XukIesjjweApNpnnUA2WR/YerWsD2P2y82yVzYfvxvGIAgAxBh33g/EAiBv8OLFC5pMJgSAUkpMRG7IAhmbODsR4bH5+a7P15h9xsxUFIU/OjqqmqbBcrlcX11d1X/5y1/89fU1r9drSinRarWiL774Ysz+uBNN0G8aAh8KQMZX4H58SN+Hn8GYfTAurtvOpv3ztp4fNgYaY14FPYwxPxYGhp4fQCL0fTqavpxVqhtwWYLqGtQ0wGwGmjR9n4+qgpQltOybnOcwHEO/j0yEhD7jYyx1lTE2XN8qeWWBD2PuBMu2vJv2JQvEAiBvcXBwABGBiBD1T8RuKHnFOWdu25aur6/x9ddf4//9v/8HItLpdIq6rlEUBchWNowB0Kcve++ZmUMIQUIIhaqGi4sLt1wu+T7cK2VZakpJx9eh7JWgD+LImBWy6/P8rm67NFYCxph386aSSiOrXbuf3tQM3cY9Y8zGpl7O7Vljxph3R0QgdiDvQXUDms6AxQFkMgUmk77RedOA6go0nUKrIehRlshFASk8svN9ySvfNzlPRBCiPqBCQ5+PocH5+ICmCuvzYcyes6yPu2lMFNjOAtk1C4B8i5wzee8p50wiwjlnHpqec9d19PLlS/o//+f/AIC2bauPHz/G6ekpee+x6/QeY/YIMTOYmZjZiYgLITgi2gQ/iqJAXde7Ps8fZOwBMgQ6VPtP6WFeffeCH6Pth3pbsDXmu7s5cR/vo+1Gfmb3toMc28GP275vjHk4dPuVXr2nv/odxpjvQ9kBQ0AD0zkwnwOzOWg2g04mQNP0fT6auu/1URZ98CP4IePDITuPzIzsHNJQ7kqINpkeAt00Nu/T84d5mT3WGGPMj0ZVNy0itqslxRgJAIUQdnZuFgB5R8OFo6HkFYsIr1Yr6roOKSW8ePFCX758qSklqqoKTdNYAMSYb0eqSttR4X/xL/7FLs/nR6GqYxksYOgJstMTMsbsle2FdAsq7ofbagvfdm0sCGLMA6evl8Gy8duYH4gI6h1yWSHPF5DFAWQ2A83moMkEmEz6cldjyau6ghShz/YIHsm5PujBjMT0WtkrUekDHkPgY/PfE30toGmMMeb+swDIW7RtS6pKzEwiQsxM6BdsWVUpxkjr9ZpijIgxoigKPH78GG3b2o5OY95iOyoM9Glxw/11rwwZIPdusWx7YVBE7OHfmO/gTeOB3Ue7d1tQygIexhjgthwPfeN3jDHfgqgPRLCDeg+t+94eulgABwfAdPYq+DGZQKoKqPt+H1IUkLHBuWOkIesjMyGpbhqdb7I+hv/k5nXT7+Nv/2MbY8xDtC8l7y0A8j2ICFQVOWd0XbcJeBwcHGC5XCKlZA/LxryD7eyP5XJJIkJ//OMf6ZtvvqFf/epXuz69H4yZd30KPykb54z5fm67d+x+2g92HYwxr1F91e+DCAqAx0wxC34Y8z0R1DmgrKBVDUynwOIAfHgEWSzAkykwnULrGto00LKElCVyWSAFP5S8csjMSIRXQQ9mCPB6n4/b//PGGGP+RnRPHrDu9+rcj+xNWR3jbmhjzA/3xRdf7PoUfnR7EvA2xuwpm0MYY8ye2wRCtA982NzOmO+PCOo9pKqhB4fQ4xPQ0THcYgE/n8PN5+D5DJjNINMpZDpFairEqkQsCrTeoXWEjglxaHSeCMhQ5CE0qbA1GmOM2RchBK2qaqeDsmWAvIMY42YBcyj3YjX9jfkRbN9H3nvNOevp6an+6le/utP3FzNbGTxjjDHGmDuOiIAbZfFsY4sxPxABcB5aVX2/j/kCWCxAsz7oQZMJZGh8LlWJHAKS7/t9dIyhyTmQFVDqe3wIABBBxqCHwgKVxhjzN7a9Xr5v6+aWAfIWq9VKY4xb/bJI0WfvWHNjY36A7UGRmZWZteu6XZ/Wj4qZQUR038tgGWOMMcbcZ98W8LCAiDHfjYIA54CyhDYTyJDpgdkMmEygTQOpa+S6QioKpKJA9K4/XN/sPA5BkE3D8+HYND2329IYY3ZmXO/bl/JXgGWAvBNmViJSVVVmluFCynZUywIhxnwvqqqac4Zzbtfn8qMZGrzT+H674bsxxpi7xRqhG2NGY+ljgmWDGPO9EaDM0BCgdQU0NWg6hUwmkMkEqaoQyxIx+D7owYTEjAhF1D7QkYfuHor+1/0vhrJXdl8aY8zOjHOlfauKYgGQb+GcU2bWnLM652QIdggRqXNOi6LQEAIODg7o8PAQk8kE3nubDBvzLYbFpDGwqN77O7+6FEIgVaWUEo2BD1W981kgtvBnjHmIbC5nzMOm269EwI2Ah77hsJHDmFsM95AyQ4sCWpbQqtwEQLSugLpCriqkskQqAtKQ8RGZkEgRQRAaMj7GSlfa9/zAGPiwz25jjNkLzKxAv66+63MBLADyTphZRUQHQkTCzBJC0LIs9fDwEKenp3j8+DEODg5QVRXu+oKnMT+VcTF9O2tKVbXrOtR1vbPz+qHath02AxIxM4nIJvhxl7NAxutlQRBjzENhu7qNMaPbZj82Phjz/QgzJARIWUGbuu/zUVfQqgTqClpVyFW5KXnVMSMSIQLI6EteieqrgOP284ndl8YYs3ecc5pS2vVpALAAyBsdHh4qAPXeKzOP2R+ZmfOQASJVVelsNsPf//3f48MPP6QPP/yQHj9+jOl0eq/K+RjzExn76dzLlXVVJSJiEeHh/a5PyRizh2xs2B9vCnxsL7BYMNiYh2eoaQqCZXkY830pM9R75KaBzBfIB4fQ2QxoGmhZQYsCKPvgRwp+yProgx99nw/tm57jluCHMeZBsPv+bhhbSOSckXMGAIjIzi+epSl8iyFVR7z32TmXnXOJmZNzLtd1nQ8PD+XDDz/Ev/k3/wb/6l/9K3r06BE1TWMZIMa8TkVEYow5xhjbto1d12VVzUQkqqree40x6s9//nP99NNPd32+38lnn31GTdNQzpmcc5RzZvTj63iMGSD2vGzMAzcusFvgYz+NNWvH98Cra2UPXcY8XJsdO0OgtB8XaNN/QIiQiSHM0LEMj43zxrxCBPEeUjeI0ynSfI40nSJVFaQqkYsCqRyCH94hDtkfiYAERYYFP4x5iG7Ox2/7ntlP+1YCy1bpv8WYAYK+6Xn23ifnXCKiXBSFTCYTPT091ffffx+PHj2i+XxORVGQbfc25hURQUpJ1ut1vLq66i4vL7vVatXFGJOIiPdeQgjaNI3+j//xPwAAz5492/FZv7unT58CALz3lFJiZiZV5eGgu1wCyxhjHoLtwMdtUzib1hljxubnY88BIgKIoczI7JCdQ2JGZsZ+tf00Zk84BykKSF0j1w2kbiBFiewDcgjIwSN5j0SMTARh6vt90BBs3PqsNsY8TLYx6W4ZgyD7wEpgvUVZlhpCUBHJ3vtERJ2qRu99572Pzrk0ZIXIdj8DY8zrVFW6rksvXrxYnZ+fX15dXV0sl8vlarWKOec0ZIcIEekvf/lLffLkif7mN7/Rs7OzXZ/6O6uqirquIxEhEWEAzMxMRA4AW1DUGENE/QLa1nBg/Sb2y81rc/N79rBlzMMzBjtujuEKBajvaxBDAEKAlCWKLiIggUQs9deYDYKCoExQ56HeQ5kB56DOQRz3mVRMEGZkychbDc7t09eYh+ttm5TMfmJmZWbtug4pJXRdBwAoy3J357Sz//Kee/z4sdZ1raoqIQQZSl91zrnWe98556JzLnnvMxGp3YjGvJmIoOu6dHl5uf7qq6+u//jHP17/5S9/WbVt26WUMhHJWBPws88+wyeffLLrU/5OPv/8cwL6DBD0wQ5mZlZVh1dlsGBZIMY8TPqGHYvb5bBsHrEfxmt185rZg5cxhoayVpuxQQEFQYgRnUMsCnQ+IDkHsbHCmE0pOCXqszicg/AQ7GBCHjKmNtkeNDQ6H/6dPueKLPhhzAN089lpnJvbXHy/jddNRCAiGHpqKwBUVbXT4dwCIG/RNI1OJhMpyzIxcwwhtM65tXNu5b1fhxCi934TBNn1+Rqzr1RVU0qyWq26ly9frr/55pvVxcXFum3bmHPOzCwhBI0x6r/8l/9Snz59qnflnlJV+vWvfw0i4q7rOOc8Bj4cAKeqbiyFtetzNcb8bb0p8GHujtsevowxD8d2A7e/CoTS0P8DhMQO0Tkk75HdVh8QYx6wsUdOYkbnHDrXl4rLPPTLGQ5xjEyMPJS8ylAI+iwrsfCHMQ/Ozfn29qaxMQhigZD9NKzjKTO/tqYXQlAAOD4+3tmgbiWw3uCzzz7Tjz76SNq2zWVZphBC55xbpZSWMcZr7/2qKIp1WZbd0CBdhtpmdhcacwsiUlUVIkpEFAEkIkohhOS9z8wsbdvq73//e/zX//pfd32638k///M/c1mW1HUdERGnlFxKyQ3lrxwAVlWGjQ/GPGg3MwpuyzAw++XmA5cx5uEZmy6rar+bffOdYXc68/B126luzDZFX9KqdR6pKBBDgDgPIe6zO4bPVt38/r8+aHg1xtx/N4MbbytNa/YbEWlfFKW36/MBLAPkrc7Pz1VVRVWTc65l5pX3/tp7f10UxbIoivUQGEl3Zbe6MbswlIlTZh7LySUAyTmXAGQiEuecTKdT/df/+l/fpXuJANDR0REVRUFENPb+cGVZ+qqqQggheO/9UBZr1+drjNmhNy2iWzr37n1bcGpP5u3GmL+xV83OXy9/NS7OjgGRmwu4xhhACcjUZ3+svcfKe0TvIcybDA9wv0dMxn9pDDJuBRztvjLm4bFm53fXuD4ushnZEULQuq71q6++2tl52WrcG3z00UeaUpKqqnJRFJGIOmZeEtG19/4qhHAdQlgVRdF67xMzy7f/qcY8aMrMGX3AI3nvo3MuhhASEWUR0Rij/uY3v9GPP/74LnzK0dnZGQGg2WxGXdc555wjIj+dTv3BwUHxwQcfVKenp9VsNivLsnRDgMQY84Dc1kh7ZH0l9scYnLot8HHbNbRrZszDoar9YiyGsaJ/Z4EPY96BEJCdQzeWiRt6ffTl4wAZylz1/9ta7CTa3HfGmIfpTaWwxvc2H787uq7Dcrnc6TlYCay3OD4+1slkkokoeu/XInItIpWq1jHGy6IoroqiWBVF0Tnn8q7P15h9xsxCRNl7H733HYCOiCIRxaqqUs5ZmqbRTz75BE+fPt316b6TJ0+e0O9//3t2zjnvvSMiT0T+4OCgPD4+bk5OTuZHR0ez4+PjyXQ6DSEEC4AY8wAR0WYHzPaC+s2MEJvE74fta/S2By9jzP23GQE2Y0L/xe2skLHJc/8tsmCIMYMxS0qGI4NAQ0XgzT91DHwM/87NLCtjzIO0XQ5rPCxr/k7RoQy+lcDad8MOdDk5Ocmz2SwCaCeTybIsy6sQwqX3/rKqqquyLJfM3IpIyjnLUDLLPq+N2TKWwPLeJ+dcZObIzNE5F4cSctl7L13X3Zn75uzsjD7//HP685//zMy8CYCoapjNZuUHH3xQ//KXv5x9+OGHs/fee6+eTCbBe29jrjEP1PYupZsL7DaZ363bghzb12VP5uzGmB3YBDoGCoD49WDHpkzPVnaIMaY3foIKbu/x0d8/ChAgOvzaVlOMMVssa/5uGa+XiMA5p957HZug75Itxr0BEeHJkyc6mUykrut0enraicjae78MIVyVZXnpnLtU1fO2bS+Wy+Xlcrm87rquFZFsD8vGvI6IhJnzEPzomLlzznUhhBhCSCEEOT4+vis3Dj158oQA8P/9v//XEZFj5jAeZVkW0+m0PDg4qA4ODsrZbFYUReGY2T6xjXngLF17v6nqa/VqRcSulzEP3NikWdD3NBibN/ed4F4Pghhj/tqtpeLGjSDDP1Rv/GZjjLnB1ln337j5edgALcyszjkFgLqud3oBrQTWm+nnn3+uAOQXv/hFvry8jKq6zjkHAJX3/pKZX8YY5y9fvvyGmeuUUpjP57PpdNqEEJjsidkYAK81QU/e+85736pqS0RdCKEriiIBkK7r9OnTp3v/qXZ2dkanp6f0i1/8go+Ojtz5+Xlg5kBEBYASQMHMRVmWfuiB7nZ9zsaY3blt15I11t4/26n2o9t6gxhjHggiYCsguhkbbmR6KNAX9iGGbsYPeww0ZtsYKBxLxtEQQNx8b3RjCcWSQYwx22xOfmcoADDza2WwTk9P9fnz5zs5IQuAvMXZ2ZkCkH/8x3/Mjx8/xunpKWKMoSiKa+/9hYi8vL6+nnzxxRf1+fm5Pzk5cT//+c8R+hXPAMuwMWaDiMQ5l4bMj1ZV1yGEVlUjgFQUhRweHt6JT7OPP/4Y//RP/0SPHz/mi4sL37ZtQUQlM5fMXKpqISI+5+xgT8DGmC1W8mo/bWqO37g+b+vZYoy551RfNWLuV2sB4r/azU7Er/qBALCpnzG3oFuCGVu3ys3NB8aYh+tNY8B2PxCzv5i5T+5T1Zz7dtlFUaiIKAD85je/2ckDlQVA3k4B4MWLFwIAR0dHGkJYhxCCql6KyIuu68q2bYu2bUMIoTo5OWlyzjPYRgVjtulQAit679fMvAKwArAmopaI0nq9zimloYQy7fP9Q8+ePeNf/OIX7vz83McYy5xzLSINgEZV65xzlXMuYEFQY8yWm5kgN/uCmP3wpkDHdpDEGPNAbAdHxx3rNGR7MIPYDV9jgPpf28KMMaPtoODN++L1gMeYa7WddalDd3TbgGDMw3Xb/Nvm5PtrLCesqnoz+2PXbHHu2+knn3wi//RP/5SfP3+eU0qRmdsQwpKZLwG8vL6+fnF9ff2ibdtzEVmpaoIFQIx5DTPnoel5G0JYEdHaObd2znUAYl3Xd6IJ+tnZGX3wwQfUdR2/fPkydF1XiEjNzI1zriGiRlVLVQ2qyrBtgMaYLbctjNli2X74tmCUlcIy5mEZG6AT86vxoW/XDBCBmfvvDQeYXmWC2LBuzGDrfvir3dsEHY7tPiC6udPGL9hnrzEPyZsCHLcFQcze0pt2fUIWAHk3CkDPzs6kLMtUVVXnnFuFEK4AXDDzeQjhPIRwFUJYO+csAGLMliGjQ5xznXNuzcxL59xyeN9WVRXbtpXVarXv2R8AgLZt2XvviCgQUSUikxjjNOc8JaJGROqUUiEiTlXtEdgYs3FbPxCze9u7S98UCLFrZszDsulZsP069PoAjxkfDHYO5IYgyKYUlo0XxrzmRlzw5h2yKS2n+iruAVtUMeYhe9vmJJuX76ex/+/wy70IfIwsAPLuFID8+3//77NzLjZNs/beX/9/9s5lN5IjS9P/OXZx94ggg6QydYMarWkUBoNUbxqafVUBs5kHyFeYfgxRL9GLeYTJbT1ACejVNBqzklaNKsyUqkqVFG9x8ZuZnTMLd4+MpJhSXUUyaR/giGC4M+hBDzc3t9/O/1trN865FRFdq+p113Xr7Xa7reu6adu2Tyml+3TAM5kfC1VVEUkhhL5t267ruialVDPzlogaImqstY0xpuu6LlZVldbr9X0/V+jZs2cUY+Su6ywAV9d1GUKYq+pCRBYppUVKqRpzQIyI5HY2k8ns2O+s896s4pvrMj8ebwqnf1NWS+7WZTKPB1X9TnizTiKHYZAxgDFga0HGAsYisUFkg0gMmYLRc/ueeeQQaNfvIWAQDLHn6b97zrvts9d/JvN42Z+YlPvjD4vx2GhKCcYYHccGVVX1d7/73Z3tVx6Y+xP54osv5MmTJ/Hp06ctEdXGmLWIrFJK13VdX11cXFyenZ1dnp2drdbrdR1CiFPQSybzmFBViTGmpmnazWazWa1Wq6Zp1imljTFma62tVbVxznUHBwdhu93K2dnZvT5XVBWXl5dcFIWJMdrValWEEKq+7xchhAMRORhFkCql5EUkh6BnMpnXMj/2H4FcEXJfmISP/ZupqSrkZkB6JpN5XEyz0HdCBhMw5n+QtYP4YS1gLdQ5ROcQnENnDAIzJHcFM4+YoR6KXlnK4ZVVHNOeW/CuEnPM/MDtkxAymczbzf690X7f+6YQkgXS+8tYBSIYRRBV1a7rsF6vcZe29zkE/U/ks88+01/+8pdps9kEAK2qOgDbpmnW33777XXXdefffvvt8smTJ/69994j772x1hpksSnzyBARCSGE9Xq9Xa1WV5vN5rLv+1Xf9xtjzBZAw8ydiPTb7TZeXV3JV199da9Hlj7//HM6OTlhAJxSsszsYowVgLmILERkZ4E1CSDZAiuTyQC3ix6q+p0qkMzdcbPMfrrpmm7AcmB9JvO42LUF+8sUhM4MGAbMIIKQdSDnINYiOA8JATEJVHuwKlg1yyCZx8de9scog+zyc3iqjtrffKwK2V1zRXL+RybzyJiEjakduHkPlYWP+wsRTQZIY/EsyfSC916LotC2be9s//Kg/J8IEeHs7EyNMSmE0KeU2hhjHULYbrfb1dnZ2eU333xz/s0331xcXFxcX11d1ev1umvbNsQYdwc/k3kbUVVNKaW+70Nd1/1ms6nH4o+r6+vry6ZprlNKG1VtrLVtSqkHEJxz8d1335XPPvvsXp8fk/1VjNF2XedijIWIVCIyZ+aDxWKxOD4+Pjg8PJzNZrPSWmuZOV+dM5lHzG3VA1OnnZkxuVvnjvzdcbP6Q0RurfbIXbhM5nGxG2TZs75SIigbqDGAdWDvQd6D3CCAqPdIziE6j2AdemMRmEc7LMp2WJnHx2RxxQQ2ZljYgJjH1/byczD0inYzv5H7R5nMY+LmZKOb5//++twvv99MlleTCHIfxsJzBcifjo6z1NN8Po9E1DNzG0KoU0rrvu+vm6a5VNV5WZZFWZZljJGXy6XO5/OCiIwxJl/FM28le7ZXoa7rervdrtfr9fV2u71smuaSiFbGmG1RFLX3vp3NZt1yuQzMnP7t3/5N/ut//a93/RHeiKrSL3/5S2rblq+urkyM0fV9X6hqycxz7/1iNpsdzmazw3fffXdxeHhYee8tM2ehOZN55NxWRfAqdDvPYroPvKn6Y7+vfg/67ZlM5kdmaKUxiCAAlBjKY+WHsyDnYIoCGBcqCkgISCFCYwJLglEBEKGiMKrYM/3JZN5+CMAofgjzUPm6t6S9TSfRQ8bH6ed89c1kHici8sZq+Vf3Upl7yM4CyxijxhgBgPl8rufn53e2U1kA+TM4PT3V09NTefLkSbq6uooxxt4518YYt9baFTNftm1b/v73v7d1XdunT5/KBx98kD744AMyxhTGmDwgmnkriTFqXdfx4uKivry8vN5sNlcppfMY47lz7gLAtTFmrapNCKHbbDahKIoEQJ4/f36v+7cvXrzgxWJhmqaxTdM4AB5A2ff9zBizWC6Xhx9++OHR+++/f/LkyZOjo6Oj+WKx8Nbat/J8zx2OTOaHuW2W0v55w8xvDNrO3B03RY/vilaZTOYxMM0+l8m+iggCHeILmGGcA1clOERQH0AxQvoeGgIkBEgM6MRBVBEBFAAKSeDcjmQeCVPvhifbK8MwxsAYAzIGwkM1iBKPlVbD9vtnyH5FSCaTeTy86f7otnuqzL1iN67HzBpjVGCoCFmv13e6Y2/lwNyPgH722Wf6f//v/xXvfSyKIohIR0S1tXbNzFchhMvr6+uL3//+95cvX768vr6+rmOM4T6U/WQyfytERFJKYbvdNtfX16uLi4urpmkuAFwYY66ccysiqo0xjbW2J6J4fX2dnj17JrjH4oeq0tOnT2mz2bAZcKrqRaRIKVUiMjfGzOfz+fzp06fzJ0+eVAcHB2VRFOZtqwDJA7WZzF/OvjCyP7iez6+7gYhgjIH3HlVVYTabwXuP/eY7V4NkMo+PXQ7Q9HxngcWANYP1lR+qPriqQFUFKitQUQDeQ5xDcm6wwrIWPRtEYkRQtsPKPA4m+ytiGGNhjAUZA7YWPAkh/F0LLIW+yv64+ZjJZB4l+/dKtGtb8v3TPUb32V/x4sWLO9mht2pg7seEiBSAdF2XUkqhLMvWOVeXZbli5usY4+Vms7m4uLi4vL6+XjVNU8cYIwC5633PZP6GSEopdl3XbLfbzWazuWrb9kpVL6uquvTer2ez2bYoijbG2BNRXC6XCYCM59R9hF68eMFnZ2cMwIQQpvDzIsZYppSqlFLFzDPv/ezg4KBaLBbFbDZz1lqTM0AymQzwXYHjtlC/7Gd7NzAzrLWYz+dYLpc4PDzEbDaDtfbWWaf5RiuTeVyoKmS3YBAveMgAGcSPElSVgwVWWe4EEHUOyVoEa9CzQU+MnhiBCNNNYW7xM287RIPt1VABYmHssEwiCBsD4mliCDCdFa+dG6MVViaTefu5rd992+SxXAlyfyEiJSKZ8j9SSqKqKiLadd2dHbAsgPxlyK9//WvZbDax67qemWsAa2PMJTNfMPOlc+7KObd2zrXGmIjcz828xRCRMnOy1nbW2q0xZmWMuSKiK1W9NsasnXN1CKEriqJn5vjy5ct7ff83XVCfPn3KAAwAZ631zFwQUamqZQihCiEUKSUnIqyqeXQsk8nsuG3AfD/cLw+o3y3MjNlshidPnuCjjz7CRx99hJOTExRF8SqI9ZYw+0wm83azH8Q8zWRXAsAMNQbqLFB4aFFAixKoKqAchBB4BzgHWANlRmKDYCwaZrTE6DFkH+TWJPN2M87WnsQP58DWgZ0HOwfYoSIEPFlgEUT3BjbHd8nnSSbzeLg5YexNfe98/3Q/GccElZmH6DQicc6piOhisbjT5jwLIH8Bp6en2nWdAIgxxs4YU1trV865S+/9uff+3Bhz4Zy7IqJVCKHu+74LIQQRSdkOK/M2MCm6IYQYQuhjjK2q1saYtTHm2hhz6b2/KIri0nu/LoqittZ2IhKWy2X6l3/5F73vF6+nT5/Sb37zG9M0jS3L0gEojDGliFRTBUiMsQwhOBExWQDJZDI3yQPn9xdmRlEUODo6wnvvvYf33nsPy+USzrnvVBGruKAAACAASURBVIBkH/JM5vEyCCE8WFcZA3UO4jy0HMSP4bGEjmHoVAxVIGotEjN6ZrRkBgGECAmUB3YzbzWDyxvtKj6MdTDeg6wFWQe2FhgFEGX+7vmg+++Vb68ymcfCzSqP6fltFliZ+8dke0VEMqIiotfX1/joo49yBchD5cMPP9Tr6+tUlmWw1rbOuQ0zX1dVdTkKIZdEdBVjvG6aZlXX9bZpmjbGGFU122FlHjwioiml1HVdX9d127ZtLSIbABtjzNpaez3lf1hrNyGE9v333++m6o9PPvnkXoeff/7553R2dsbL5ZKdcxaAExGfUiqIaBJBypSSTynZXAGSyWTexNRRvy1YO3fg7w4igrUWs9kMh4eHODw8RFEUMMbcGmCfb7gymccDTTkd+3kdzIBhwFqIc9CigBQeKAugLEBlAR0tsOAcxBgkw4jMCDxaYNGYA3K3Hy+T+ZszZHyYQfxwDtZ5WOfBzoKsHc4lfhWCLgBENUd+ZDKPlH1b4Ju5H/uPmfsJEel4/ERV1RijqqpFUejBwcGdtuz2Lv/4W4Isl8vUtm04Pj6GiKi1VkWEvfcFgHnf97PLy8uZqpZ1XePo6CgdHx8vZ7MZMbO56w+QyfwliEhq27a/vLyst9vtar1eX9V1fR1jvGbmaVkZY9ZlWdYxxm6z2cTlcpmePXsmP//5z+999/abb76hg4MDw8w2hOABFABKVS1UtRARH2PM1R+ZTOZW3hSeTUQQkdyRv4fsV3rsCx831+Vjl8k8DnZtNxFUgQRADEOcQVIL9g7kHeA81A8ZIPAe0nUQY6DGgChCMWaIILcdmccADfZX1oKdBZwD+2GBdRBrhmoqZigTBAoZItAh+/Kg6isBMpPJvPWoKpj51nuoN91XZe4Pkw0WxmIQY4yoql5dXWGxWOD58+d3cuByBchfhp6enuqXX36ZAMTtdtt775uiKLbW2rX3/toYcxVCuLi6unr59ddff/P73//+5cXFxUVd19tuSFCPIiLZDivzkBgr2iSllEIIoWmadrVarc7Pz68uLi4uttvtpYhcee+vAaxijBsAWxFpAfSz2Ww/++Nef/e//PJLOjg4IGY21loLwAEoVLW01pZFUZRlWRZFUXhrrcPQruYeeiaT2XGzjPumt+1t22bujtuqPm6+lo9TJvPImNpxDAOzyoREBLEWyRoka5Gcg3gHKRy02KsAsRbCjMQEYR5muNM97wBnMn8uU7XUmJUDM1R6sPcwRQH2frfsMkAMQwmDvRzGG0RV7KLP8zU3k3k03FZpfXMCWeZeoaMrjIQQpO97iTFKSklERJh5F4B+eHiofd/fWfcnV4D85eiLFy/kk08+0X/6p3+Sd999N3355Zd6fX3NROSdc2Xf97brOg4hEACy1qKqKkNEaSwFKowx1hiTq0EyDwJVlRhjijGG7XZbbzab9Xq9Pl+tVt9uNpuX1tpvrbXn1tpL59wKwKZt28Za23nvw9dff51+9rOfCRHd+3u/58+f4+uvv6YnT54YEXFjxUdpjKmqqppXVTV3zs2fPn06Ozg4KLz3hpnfmqty9tfMZP467Ftd7Zd0Z1ul+8ckdojId8rwgZwDksk8VhQATUIoEYSApDQM4FoLcg7wDuo9xHukwiO1gwCi0yx3wiCc4AHMAspk/hyIoMxD5VNZQsoSVM1gyhIoS3BRgooC6ocwdFg7nhu8J3zshR/f9efJZDJ3wtT3FpHdzzf755m7R0SQUpKu61Lf913btl1d130IIYpICiHoJICISLbAegvQ09NTnJ6eyk9/+lNst9s4m8167/2267prEbExRmZm9H3Pq9UK33zzDfq+709OTmS5XB5WVVVlASTzUEgpSdu23WazqTebzfV2u71q2/alqp45514aY14WRXHOzFfOuY1zrlkul31RFPH8/Fx+9rOfTfd9956vvvqK/uEf/oGJyIQQvKoWzFx672fz+Xx+eHi4ODo6Ojg6Opq/88475Ww2s8aYt3IUMw/6ZTJ/OjfPmdvOoduC/jJ3x27Q5RbxA8gVIJnMo2VqG4ggqkhEw8T0MeiZmEDWAN5DiwLqCyTnkEbxA+MiewJIJvO2oVNlVFlC5gvowSFoPgdVM1BRgAq/s4hTN4iDYAPwq/NLASCLH5nMo+XmPVEWPe4vqqpd16Wrq6t2tVptt9vttu/7pm3b2HWdWGunahA9OjrSly9f3tm+ZgHkr8dOBPnggw+SMaZPKTWqunbOMTD4oKWU+OrqCm3bou/7NGaFGGY2zGzHmeNE+c46c88YbdpUVXW0vWqur6+v1+v1xXa7PY8x/oGZz8qyfMnMZ8aYC2vtNTNvvffdfD6PH330Ufq3f/s3+fTTT/UhVH8AwE9/+lOcnZ3RZrOxqurGwPOKmWfz+Xz+/vvvzz/44IPFwcHBbD6fF2VZvlUVIJlM5q/Dmy7rtwWjZ+6W6eZKRF674botuD4ft0zmkTEOziqGoOY0Pmcesg7IWsBawBeQooA6B7UWMlr9yCSA7N5nCH7etSJ5cCfzUNizq9pHjIFYh1jOoIsD4OAQPJuDqwpUTtUfo0WcdVBrhvNh6g/tzfbO1leZzONkfzIS8ObqjyyI3D3j+GBcr9fdN99806zX6zrG2FlrgzEmMbOIiFZVpaqqz549yxZYbwl6enqK//W//pcsFov4m9/8pp/NZvVY/UFd1yGEYGKMtN1uiYhQFIWdzWZ2unn23vtsh5W5j4iIpJRSjDHWdb3dbrer7XZ7ud1uz5umOWPmM2Y+s9aeG2MunHPX3vt113VNjLH/6KOP4osXL+T58+cPwvpq4uzsjH/729/aoihcjLEQkVJEKmPMzDk3m8/ns+Pj43K0v7JERMw5XimTybyZm+F9eRD9/rAvftysArntOOXjlsk8TqYwcxoHaZVGAcSYPSssB/EeMoogw0x3RmJGIkIghoWAVXcBcrlFyTwUhjycYRmqNobsDzEW6jxSWUHLCjSbwcwqUFmAy1fihzqLZBmyC0AHksiu0iqLH5nM4+Q2UeNNokfuh989qqoxRmmaJqzX6+7y8rITkb4oilRVlTCzWms1hCBnZ2f4f//v/+EXv/jFnexrHqX766PPnz+X//2//3c6Pj7uF4tFU5bl1lq7KoriyhhzrqovU0rfNE3z+8vLy9/94Q9/+N0f/vCHP5yfn583TdOklOJdf4hM5iYppVTXdXd5ebk+Pz+/vLq6Oqvr+mVK6SURvWTml977M+/9t0VRXFprV6paW2u7s7Ozhyh+0OnpKX/99ddmNpvZlJIHUKSUqhDCXETmIjIjotIY46y1bIzhqYrrrnc+k8ncH25mfQC5836f2Rc8pioQ4PvD6zOZzONhP5cgjYswDSKHHYSPyQKLigKYBJBRBBFmRGPRMqNlRkeMiGyJlXlYKIAIQkeMhg221mHrC9S+RFtWCEUBKUtgrPigshxsr7yHuKEqSoyBMO0qQEDZbjeTyeA7lR837a9uey1zp+jehOkUY0wiMnWRkrVWRERjjAoAn3322Z0cuFwB8jeAiPT09FS++uqr9Omnn/YHBwfU9z1ZazHmCBAATinR9fU1N02jdV3Htm3Fe2+ttcY5Z/HKCivfZWfugtF+dXgYba/q8/Pz681mc9627ZmIfKuq3xZFcWaM+ZaZL6y1V865NRFt5/N5IyL9crmML168eDC2VxjEDwLARVGYGKMF4AAUACpjzJyI5kQ0U1WvqtPEvUwmk7mVfeFjP/A8V4zdP/bFj/2fv2/7LIhkMo+IPRssGgduhWjI+DAMtm6oAikKwHuQ94MIYgzMKIREFfRqwAlgUhjkgd/Mw0IAJBoEkMAW0Rioc0PIuS9gnId3DnBudw5MuR/JGiQeqj+EeagkmYRFomwFl8k8cm5aYAGv+tvMDGbe3U/lPvj9gYh0tLwSZk4iIsYYiTFKSkk//PBD/eCDD7IF1tvGZ599pi9evEhN02C5XFJVVdQ0DQCYlBI555BS0u12i+12K0Qkxhgsl0tnrVUA6r13xhjHzPk4Ze6EfRV3sr3abDYXm83mPIRw5pw7c86dGWPOp9Bz7/21qm4Xi0WzXC67L7/8MgKQ09NTuevP80eyEz9OTk7MbDazdV3vxI+qqubW2sOqqo6Wy+VhVVUza63NuT2ZTOaP5bYybsqzHu8N+2JVSulWAeRmKHomk3l8TG0DEwHEUGawc0BMY85BNzy6QRAh50EhANZCUkI0iqAKpzoO/ua2JPOwEBAiMwIzgjFQY8HWgsfvvDoPtQ5wowDiHGQUAZMxiERDBRUNFlh5Rncmk5nYbw+ICM45zOdzWGtxdHS0e56HYe4HRKREpKqqRCREJNbalFISa60sFgtNKekvf/lL/OxnP7uTfcwD638jxgMvL168QEqJAFBVVbi+viZrrYpIDCGklJLEGGW73WpRFHp5eWlUNaWU0nw+P6iqap4FkMxdMA78pKZp+qZpms1mc71ery/rur4IIXwrImfGmG+MMd967y+stRfMvHbObbz3TUqpvb6+DgDSF1988VDED0zix7Nnz7iqKnN2duYAFE3TVEVRzGez2eHJycnRwcHBO8fHx8eHh4cL55zLAkgmk7mNP6Zp2A/Tzk3J/eBNJff763MIeibzuFEM5b8iowjCBjB2EDuSAEUB8gW4KCBuqASh0AMhDMHPKsPsd5EhPwGEbISVeSgoCEqDCJKIEdnsqpzgHNQ5iLNDHs5Y/SHWQqxBZB7Ej2nB8M3XXP2RyTxqblpfTc/H/GQsl0vM53OcnJzg6OgIRVHkfvg9YHR6USKSqQIEQBorQURENKWkv/nNb+50P/PA+t+QPREkAtCqqsQ5J03ThK7rOgBBVZMxRlRVt9ut/Pa3v0XTNKFpmvT++++Tc66wNh+mzJ2gMcbUNE3z7bffrkfx4zyE8C0RnTnnXhpj/jCbzb6dz+cX3vtVjLFOKbV93/fPnj3rAaSf/OQn8vOf//yh9GTpyy+/pE8++YQBmKZpXNd1XlULVS2Zeb5YLA7ff//9d54+ffpkPp8/qapqXhSF40fgY5NnZGUyfx438z9uywHJ3B/eJH6IyG6mWZ6lmslkgFc2WCACDANqQOpBikEAKYvBEqgsoV0Hdh7sApASVGRYaBhI3r1hJvMQoDH8nGjI8WAGjIHsrN6Gyg91Qy6OjI/JDPZXiQkRQ/WHYm/AM4sgmcyj5WZF/GRH65zDbDbD06dP8eTJE5ycnGCxWGA2m2U74XvAVP2BQQRJk/0VhihhERE9Pz/Xjz/+WD/++ONsgfW2Mn4J5Pnz5/hv/+2/6fHxsc7n82StDU3TCDCc1KqqXdfFEEIE0AHoFotFdM4FETkUEQPAGGOMtdYZYywRmTzrPPOXoqq7wCIRiVNDpaqx67p6u92u1+v15Waz+bbrunNmPjPGnFlrXxZFceacu7DWXnddV89ms/b8/LyvqioCiET0YCo/gKH643e/+x0DsJeXl46Zy5TSvOu6g5TSgaoeENHhbDY7nM/nhwcHB3NrbcnM/Dafi3mQ7wGzH7QNDDeVu1XfPa53/TV+fZf2fngLTq+b/9vJw3bsA9z5/z7zipvix5sssParQDKZzOOEQAApaBqAMWacyq6gYqj+QFlCyxLoeyBGUIowqoAOAghSAoSy+JF5YIyh5aPwQdYC46LWjnkfbgxBL6BFMQafWyRmRIzpuKqIow0cgCx+ZDKZ1/rgIgLnHKy1ODg4wMnJCU5OTuC9hzEmCyD3BGYWZk6j/VVi5l0IujEmee8lxqgvXrzA8+fP72QfswDy46AvXryQTz75RP/zf/7P2jSNMHOKMTIRmb7vjarSGAyTrLXBOdevVqtIRE3TNMuUUkFEhXOums/ns7IsZ9bat3rQNfPjoIPnWmyapmvbtkspdUTUE1Hb9/22ruvrrusuuq47jzFeOOfOAZwbY86Z+co5t14ul1vnXNu2bQAQvvzyS3n27NlD671O1R+mLEu3Wq2KsixnMcZFjPGg7/vDEMKBiCwAzKy1pbXW27e8ROtmTkHmATDOnrv14iCyW3fr+v2guT/yz/0xl6E/6vuje5URUEyf4DVP9Glm4ANnf4B9P8AvX9LvD/tB6DdFqv3jltvGTOZxo6N5lU6z4ZkBO7QNXBRAUYDLAigLUF/uBBASAUIAWQFSBNIbr8yZzP2FCGAahD9jADtawI15H/BjFYh3SLvsD0YiQtSh+iOJDhVQY+VHvqpmMo+X/ar5qfpj/57Je4+yLFFVVRY+7glT5QczyyR+jBOhU0pJjDGSUtIYo/Z9r+Pv3Mm+vtUDd/cMPT09xenpqfz0pz9F0zSYz+fddrs1IsI6nOmBiHoRaeq63p6dnW03m80lMy9DCHNjzMFisTh677333hkKQawFkM/6zF+EqmoIIa7X6/r6+nrdtu1GVWtjzAbAquu665TSlTHmgogumfnaWns5/rzuuq6u67oriiJst9v06aefyi9+8YupBO5BcXx8zPP53BCRs9aWIYRF13WHKaWjGOMyhHAYQpillLyqch6szNxHvlNpgHHAdnpBB3GBbm60h+ofOwyj3+tYvnP0UMX3vePudldfeaoDe4PMuzekV/YID4ibGR/7S67+uL9MAsht1R/7Nlj5+GUyj5ddeyACZQDEEBIYNVBrQd7DlBW07MAhAimBUoImGcQQSQDzMIj8oOqmM4+eSbRgBgyDrAHcqwB0+CH3Q72Der8XfM6j9RUQoUP+hwKi4wnwAPt5mUzmr8MkfEx97+n5NCFpEkUy9w9VVWYWY0wSkV2RX4xR+r6Xk5MTaZpGnz9/rrijmtcsgPy4vCaCbDab2HVdZ63lEIKKSMJgG9T1fd+uVqumrusNgGUI4cB7f5hSahaLRSyKIhLRgoic6tDdVlWaKkJUh3kU4yMAEBGRMYastcYYQ0SUxZNHxGR1JSJJRJKqCgBNKcW2beumaa632+3VdrtdicjaOXdNRCtVvR4rPa5EZMXMa+/9ylq7Kopi65xrV6tVmM1m6Sc/+Un6/PPP9fT09MGJH8+fP+d//Md/5LquLRH5vu9nzHyQUlr2fX8UQliGEA76vp+HEAoRMXvnVyZzZ6iO4avAK9uNQfUAVDFcIF5tP4kLU7UH7a14NcP9zX/v1WDvK6uCHxJAhs0Et4kgOv1BIugohUzvR0y7fSHmV5ZDe5/9od0k38wDAYAYI+q6xtXVFYwxWCwW8N7v8iYyPx5EBGstyrLEwcEBYoyIMe6Oxf7xyFU7mUxmd70CxusYoGwgDBg3CCBUeJjZDJTSYHcVIxAjJAZQDIM1FuUKkMxDY8q+GeyvhsoPDy4KUFGAvB8FEI9kLchZJGsghgcLLFUIAaIKJX7V/8vX1Uzm0bNfLb8vfuQMvvsJEelogRWJKBJRApCcc4mIUt/3EkLQ9Xp9Z+IHkAWQu2AngnzwwQfx+PgYALQoirjZbIIxphORJoRQp5S2RLROKS1F5MA5t2Tm7Wq1aowxdQhhAaAQEauqRlV5HJTlMTOE98QRds6ZsizNYrHwRVFYa20WQB4RIiIxxti2bdv3fRdjDMwch/iZblvX9VXTNFdt216JyHVK6YqZr40xKyJaOedWADbMvHXO1d77LTM3McbeWht+8pOfJAzf7ztt1P5cPvnkE7q4uDCLxcKFEEpVnYUQDlNKxzHGk5TScd/3yxDCPMZYjOdc7qFn7pT9yo5R/QapgichRGUoExQZLKYmMWESSYBX1SD732b6IS9y/Z6f9vbne/b79d8jCBS6s8ACwAzVYWahAoNP+mjflfZEhCk48yEORE+znLquw8XFJYwx6Psex8fHODk5QVmWcM7d9W4+KogIzjkcHR2h6zp471HXNfq+39147ZfcZxusTCYDYLxmjSI+AWp4sAMqPMysAouARECqUEmQFMGhB4cAMi1AnPWPzMOCADCD3CB+sPfgqgQXBUxVgcsSVJYQ58DeQaxFshaReaz8IAiGwqep+iNfTzOZx8u+7RXwXTva26qyM/eDKf9jXCIR7SpAQghSVZWs12s5Ozu70wOYBZC7YRJBEgB473U+n6eiKGLf96Esy56IOgBdjLFzztUxxo0xZhtjrK+urjYxxgtjzIGIlCklLyJeVV1KyQOwImJFxAIwAIyq8mw284eHhwUzkzGG3/LogswNRET6vu/X6/VmtVqtu66rjTEdgBbAum3bFRFde++vAVw7566IaGWMWQNYM/MGQAOgYeZ2zAjpf/WrX8Xnz59HAA/S9goYKqZevHjBv/71r81ms/EASmvtLKV02Pf9cYzxOISwtNYe9H0/izH6UWTMZO6MSfwYy/2GBaMvoiSwDK8ZVUAEJKNYMr5ONP3u8CY8vQDslIk3iwqvV33cPPHpludys8M62l0pMIgfICgNftCvLBXM8HvGjNsN25tR+Li9puR+ctv/cho8b5oWL1++xGq1wvX1NT788EN47+GcywLIjwwzoyxLPHnyBN57HB4e4vLyEufn52iaBimlByu4ZTKZvz5TJeJkB6nMQwEmA8IMHkOgX4WfC2QUPlLbgVwPtg5DYX5uVzIPCCKADdgOtldaFDBlCS4HEYTKEjpWQIm1UOcG8YNoqPzAMKFlV9V7l58lk8ncOfvixr74kVLaLVkEub+MGSCvBZ+nlMR7L0VR7Ntf3Rl5BPzu2BdB9NmzZ/Kf/tN/Sr/61a/SYrGIAIKIhJRSn1JqnHO1qm5EZNO27XXf9wfMPE8pVSGEmaoWqlqklAoAHsBODJmWrusKAOVyuUze+9IY40fbrMkya/e4/9rIbT3y77xGI8aYXS9eRCSl9J2qgD919vwfGbR753cO3ycC/DGN9c3fJyLigekYiYiIDux+Z//53nsME9GINITQ931f13V9tdlsruu6XhtjamNMDWCtqitVXXvvV0S0YubrsizXqrp1zm1DCI21tq2qqluv1+HJkyf9H/7wh8HCdQg5epBM4gcA45xzIuK7riv7vp+LyAGApXPuuCiKo8VicXh4eDgvisITkUG+U83cITuzjEkIUYUBgVICq4KTgCSBk4BVQGmYeboTQAAQpkfC2MS8stP63j/++jb7jdZ+7sfNdxpEEN3ZWsl44ysYZswKCMLDDbUaBkRgrB22YQbxOFMQtBNtdsLKA7DDum3gXFURY0DbtthsNgAUs9kc77/fIaV0Nzv6iGFmOOcwn89hrYUxBiEErNdrdN1wTPatr/JNWCbzuKH9ykXsOt4QIrAxUGuAwoNFxioQBXcdtO+HGfJtC1gzZIDc82tYJvMaRCBmkLVg54GyhC0rcFWBqkEIQeGhzkGdQ2KGGIOkMuR+7FVQTtW8mUzm8XKzqnqypTXGYDabYT6foygKGJPnod4zpjFHMcZEY0y01kaM+R9EJDFG/fu///vd2ORd7WgWQO6WyS5ITk9P+enTp3JxcSEikg4ODuJsNgvM3Pd933Rdt1XViohWdV3PY4xzEalUdRZjnKtqJSIlgGkpRKRgZqeqnpktERVFUVR1Xffe+xJAAYBEZJchgt1k4lfCyPT6nuXDbj3wKm8EAJiZrbWmKAo3Zoxo3/ex7/uUUtoNku///hv/OXtixo3Bhjf+4p8jgNy2H39JB+y2E3p67aaqfdu2+68TEVlryXvvrLWGiKbMjjjmeEwNyJ5tKsn0GhGJqgoRpdH9qm7b9rJt28u6rlfMvDHGbCZ7K+fcmog2xph1VVUr7/1WRBrvfQug22w2oW3bsFwu43/8x3+kL774Qk5PTx+s+AEAn3/+Of30pz+lr776yqSUrKp6AKWIzFNKB8y8LIri6ODgYHl0dHT49OnT+Ww2K8bjke9UM3fDvvUV0TCgogBLGh5jAqfXF0oJlAQ8ZYOM7RFjEBJozADhPfurW7/ge1/7783+oD0RRF/d3E45HyLj81HESETDzNnxBhnWQGWcGWgMErCbIUtMw83za3+PHszswd0N/zi7KSVB27ZIKcF7j6apEWP83iyWzN8Oay2stXDOIcaIqqp2GSC3WWABeeAmk3nsKMbBm+laxAxlAZwbAtJFBwssEaArga4b8kGcAxkDNiZPq8k8KAgEMgy2DlwUgC9gqhJcVeDZDChLaDFUgaQx/yNOk13wahLMLgsuk8k8Sm7rQ0+TxoqigHMOBwcHOD4+fq1Pnrk/jBkgaRQ/QoxxZ4HV973UdS1N09x5Q58FkHvC6empqKqenZ3p5eWlPHnyJL7zzjv95eVlJyL1bDZzKSW/3W5LVS2LoihFpCSimarOU0oVEVUppcoYU4lIxcyliBREVBCRK8vSAyjW6/UspeS9937MDDEAWEQMDaUEPC0YBRF6VZc9Ba2/JpaM21NRFLYsS79cLufOOSMiWK1W7Waz6fq+D5OgMokrN8JEX2vF9qtS/lwB5Icaxu9b/0ODGW9a/0MCyI3qDBCRTl6He+sVAKy1VFWVPTg4KGezmQeAtm3b1WpVt20bUkpp3H6qwhBmTqMIkpg5AohE1ItIG0KoY4wra+11WZZrY8yKmdfW2msi2nrvN6q6BVAD2Khqy8z9yclJ+Prrr9PV1VU6ODhI/+f//B/56quv9KGLH6pKn3/+OTdNY/q+t6OVXAlgJiKLEMJyPp8fHRwcHH/88ccn77333vG77757eHh4WMxmMzNV5WQyPzZEtAs5JwV4tLriJLAioBhhQgSnBBMjKASYfREEgwDCOlSB8Ch8DC5Yr9pbmv4Wbhc9vi/7Q7FXATK0gMPNrg7rRAQCRcJY1cEM4SEYU60FnAPckPshGPYvAYAhJJFhEFpfD01/CNyc2XSTG1fCv/0OZf5k9it5svCRyWQA7KoQVYfrGgNIhsFqYL0fNoEOeVZdD2r7IS+hLgabLOZcAZJ5WBCBzZD/YcoSZj6Dnc3B8xloNoNWFaQsIKMFVmRGZEZShUga7E/H/uFkJZfJZB4fu/vO8Ro6jY1ZazGbzfDkyRM8efIER0dHODw8RFEUGKbb0QAAIABJREFUWQC5ZxDRNA4ZjTHBGBMGI6DBAqvrOl2v13dumZ8FkHvEaGMkn3/+uf6P//E/0i9/+ct0eXkZnz592p2dnVnnnF0sFnVKyRNRgaHKowIwU9UKQKWqFTNXqlqNA7k7AcQY4wH4tm19SskxsxMRS0RmzAuZhA+z95yZmW57xJ4gMlWRlGXpVLWYz+cLADalhKZp6s1m09Z1HYGdoPGa9dYtlltQVeIhUHBfG/lB8WO/MZx+/7btbm57y/t937qbNlVv2vjm6zfHDnUSPfbFDxEBEan3nlJKzlo7s9Z6ItKmadrNZrNp27YLISRm3uXHjaJHApCIKBFRABCIqCOiVlUbEdmOFR5rZl5Za9fMvDbGbJm5jjE2zNx47xsi6ufzeTw5OUknJyfy4sUL/eKLL/Szzz6788brr8Hnn39Oz54941//+teuLEuvqmUIYWaMWVRVdVBV1XK5XB6dnJwcvfvuu4cffPDB/Pj4uCqKwlhrOV94M3fCOPiqOgoXOs4qjQlmFD+4D6A+gGMA+h4cIihGIMZX26uAdQiKYh0qQ3iyxKJhhvt+lcnN5vf7qj+GG9m931DdWVWp6mB5pYo0bpPGvI9pSaMAQkUJEQF7D6iDGgMzZYSMmSWT3cg0g3BUlv86/+u/MtNxuyH+76pv7uluP2puCh253c9kMreyV4U45YEIADUMhYWIDBUfMQGFB5UFqKxAZQEUJcQXkBAgKe3C0vOs+MydM17zpgw2HftfxIzkHaTw4LIaqj3KEmZWgWYzUFUhlQXUD+JHMgaJGRFD7sf0fkM/Ll9XM5nMq8p4AMP9H/Muj++dd97B8fExnHPIWcb3i70J3MkYE4goTEHoxpgUY9QYo37xxRd3vatZALlvTF+e09NTYOhrAABUlf/n//yf5vj42H744YeWmV3Xdd57XxNR3XVdCaDsuq5i5oqISlUtABQppYKInKo6VbVN09i2bW2M0TGzwfA9MGMFCGMMTZ+W8TVmZiKiXWXICE8WWKMQ4owxRdd1i5SSFRHUdd1sNptuu93GVx9zN4LwmrXW+Fn3xsxes9d6o1Cy/y+cnty0qLjlfV/bZp9Jdb6Nm9ZVtwkBk4Cxv83UoO9Vg+wqQfbW7yytVFWdcwTAzWazqus6T0Tatm1b1/WmruudAKKqsi98YCg3i8w8NUAtEXXGmJaZG2vt1jm3BbApimJNRBtVbZ1zjaq2RNQxc/fxxx/fmvExfj/fBvjy8tIWReHbtq1SSjMimjvnDpxzy9lsdnR8fHx8cnJy9PTp08Xx8XF1eHjob1YrZTI/GjtLqb1A89FSg1MC+gAKg/iBrgP6Hug6aAjQEEApQVMCRPYqSBQcI0wMMCrYlz6+TwAB3lwBcpsAsrPAmnI/VEDMgLWQUfBQa6HGgJyHOAfEBJIESWkIdvd+EDuMGW7CDb8Wjr4fRHtf2RdBXl9eXef2qx4zd8v+sdr/+aaQlclkMhPT9Y4ACBGSGXISKAnIJ1BRgKtyyEmoZkA1g8yaIfdJBNz3MJIGESSTuWMEo4/JWKkLY0DGQMsKOpuBqhI02l7xbMj/QFUCRTFkfxiDxDQs43vtBBXkSspMJoNb+9U0ZoDMZjMcHBzg4ODgjvYu80MwsxhjEjNHZg7MHFNKiZnFWivWWnn27NmdN/ZZAHk46PHxsQBIzIyzszMURYG6ruG9V2ttTCn1ItIRUc3MXlW9iDhmdkRkU0oWgCEiq6rGGDPZXxkac7ZTSmZSOkSEmXlXBULDKD2Pg7+TiEGjDRCJCKeUTAjBbrfbwhhjRAQhhAAgGmMEO6t2ek3YmAQJESFjzHfsryahQlVpCj0Ske/8PjO/9vrun/fdzJIdt4kgbxJAbnudmW+zvHpNAGHmfZur14SPUd1WEZnW7UQQYwxSSqZtWzvmuEjXdSGl1I3/0wRAJxFkFCp2IoiqRlWNzNwB6FW1V9WOiFoRab33tYjUzrkGQKeqvTGmX61WMYSQPv7449244lsIYRBA3HK5rERkrqoHIrIsiuL45OTk5P3333/yzjvvnBweHh4dHR2VRVHkNjNzd+x3DKf8DgIgMggbXQd0PaTrgLYDdx1i2wJtC+p78CiAmGn7aZZNCKC2gW0bUOgHf/Kbf/pPmJ33ennc/otTWPvola4KdRZaFEjVDKEskHyJaAzgPeA9qOuBvgdVFSRG6Bjkzs6PN8wWsldBsfvbD8xKYX+APYsf95O9SQwAXg9qzIM3mUzmJlNbIaqDCMIMMsPgsXEO6ofKD8znkK5DiBFKDCGCwwbU9zDfMyErk/mxECIEInRskLyDeg9TlqDZAjg4hM4X4PkcNKtAo6CnZQn1DuIMxBokorHy41UWHPD23mRmMpk/npv96KnPLSIYx8hyX/ses18BMk6+DqMTTSrLMvV9L8fHx/rFF1/c+UHMg3kPiOfPnyuA9OLFCwBA13XqnJPZbBa7rgvjDP+GiGzf946IrLXWxBgnwYNFhFXV8AiG7I9dlcf4SKrKxhga1+3yPiaxY2IUG15bQgi83W4NBvtb9H0vIgJjjE6/M85y3RdDML2OvUnD07rbRA5mxr4YMgkZk4gyPb/5+ze4dZTJGHOr2PGm18d93Z3Q1lrd346GUKBpnzDoSqoiAufcTgiZBJBJVBmFEWqahmKMpKqaUkoxxknk0LFqRJhZpkdV3QkhIpIABFWNRBRGT74eQI9R9Oj7vmfmsN1u44cffhh++9vfps1mI59++ulbYXV1k9PTUwbA8/nc9X1f9n0/6/v+QESOUkonxpiT2Wz2ztOnT0/efffdo8PDw4W11jrnHq3tVe503CP2wssxBarGCPQ9tG2AukFqWkjdgLpBAEE3CCJTDginIWBbRKB9B9Q1sF2Dug5I6a+zn7R3Y6vfWTUs3g03y4sFtKqQihLJeagfFq76oaIlRiAlqEyffbTA4qE8WjAKB9ibof/X+RR/E/YH02kn4Lyu2WQh5O65TeAY+zM5BySTyXwvu9nt48DvWOYHWAPyDlwWMPMZNAZojLttVAQ2BCBFIP7QX8lk/rYMVbaEyAadMQiuAKoKdj4HLw5gDg9hDg5A8xl4NgPNKmhVDpNb3GB9JcwYZ+bt7K8kXzczmcwt7FtgZeHj/qIjIiIxxhBCmCbjt8zcEVEoyzKGEMR7fy8C0IEsgDwYJoskjMNIl5eX+nd/93dydHSUuq6LxpiQUjIiYrz3HEIwqmpEhK21nFLiYYybiZkpxshjhgFZa2moTmIyxlBKaSd8jMICOecoxkjj9tM+vSaGTJUbfd9T3/e7FQBgjNlVfIzPX1u/bylERJRSmrYF8F1RwzmHm7+HW4STm8+n97353j/0/08/MCB4owrkOyf3tD4Ns653FljGmN3zUdzAzddEBNvtVqftdSjJEWPMTkgZRY/dc2aWCWtt8t5HZk4xxgQgiUhk5hhjDNba2DRNWq/XqSiKdHl5maqqkv/+3/+7vIXiB52enhIAPj8/N0VR+KIoShGZi8hh3/fLlNIRgCNmXs5ms4ODg4P5YrGo7nrH7wO5A3K3vFYhMFprDBUVMlhFhQBtW1DTAnUN3daQphlea1to14LjICYYEbAIWBKo74F6C9psgL4D/bUEkD/mMzkH7jrYFBG7HrHsod4jeg8tS3BM4CmvZFIIrIEyA8xgHkQPNgyZbMH28kDucxXITRulSfAY5hlk7gv73Yz9NjCLH5lM5ntRhRJBFBBiADLYNBoD4zzURaAsR4FfBqvHFEGhg27X0DZfCzL3Ax0rmIK1Q//Ml0A1h50vwLM5aD4fxI+qgpYlpCgg3kOtgYzZH6+JH9Dd+ZGvoZlMZron2nNMeU38yO3E/WMcu5Su60Lbtl3TNE3f983oVNNba4OqJmOMhBC0KIq73mUAWQB5UNCr7IjJlkj+/d//na+urqSqqti2LTdNw0VR0Gw2467r2BhDxhjq+54m4WESNLquI2MMqSo554iZd9s556jve/LeUwiBiAjTc2ZGURQIIdA4CE8hBPLeY1y/EzW894gx7tYBgPceREQxxlvFDwCY1k1CR4yR3vR82u6Hno//u9fed/89vo83ZYVMWGv3nFe+20JbazWEAGMMQgi77SfRYnpeFIXur5+ej0LIbjvnnIrsNI/XfhYRtdaKiGiMUZxzMimvU2VI27bivU9VVaWmaeSdd96RqqrkX//1X/X4+Fi++uor/fnPf/62XWno9PSUPvjgA7Pdbu3f/d3f2dVqVTZNM2fmwxDCMsZ4nFI6CSEchRAOUkqFiJi73vH7SO6I3B2vhA8dsjySgFIE+gC0PaRpQW0HbRpoXe8EEG5q2K5DFXu4lAbxQwQmJXDXDZUWP/JxNSJwXQcFQfshsD0UQ5CmiAwVH1MlhDFgY0HeA8YCNgKGx6pAHUpiboSL3/dv6avL3/4jvWavlLlbbjsOuyqjPDMtk8m8ial9nypAmMDGDB4R1oILD0gC0jCJASGAuhbsyyFjgb7/3iOT+dEYpjwCxgDWgosCXJbDMgofVE1B6IP4kZxFZEYkQqShimSq/FDK2R+ZTOYVU1uw37e+KX7k9uJ+ISLSdV24urrarlar6+12e9l13brv+5qGPOEgIskYI23baghBP/vsM73rLOEsgDxA6FVINv3iF7/QZ8+eyWazwdOnT+l3v/sdffrpp/jVr35Fi8WCRqsGWiwWODs7240MVVVFAGCtJVUFM9NqtSLnHKWU4Jwjay2steS9x3a7JWstAUBRFFgul9hsNt95PxGhxWKBpmnIGEPz+RwA0DQNHR0dAQBmsxmapqG2bXeCzN77oG1bmhTCruuoqqrvPAeAsizRdd0PVn2UZYm+778jchRFcevrfy7ee+267tZ1bduiKAqoqnrv4b3X8bXdY9M0KIpCj46OtK7r3T6qqpZlqXVdY3oUEZ3P5ztRJKWkRLR7LaWkKSU1xmiMUZfLpcQYFYD2fa9Pnz6Vvu+1aRpdr9f66aefKgB98eIF/vmf/3mq2n+rmCo/vPem6zq33W4LAJUxZpFSOlTVI2vtsTHmxHt/ZK09VNVSh5ycTObOUbzu2aeqMAqwYhhACWFY+kEE0TH/Q9sWWtegpobrWviugQ8BZnDcA4sCkyDyI3cuSQQmBBSqQIyQsToFKkgYNQ1jwGygzkGdB7wbwmSthVgDYgYxgUA7e7Cdn9Q97SzvV33sv5arP+4XP1T9MT3PN2WZTOZNKHS0hCQIE6IQ2Fmo+sG+MQkoRnAIQNNAiwLqPcQ5UG8B6C5Ha+qdT/L+3gyvH/1zZR4XRAQecznJGrD3gxAyhp+jHASQ5Ebxw9oh94OmEHV9Xfy46w+UyWTuDTeFj2nZt8HKtsD3CxHREEJYr9f1t99+u76+vl4B2BpjWmttx8zBGBO7rpO+7/W//Jf/ci+a/SyAPGD2wmb+IqaqiM8//5w+++wzvHjxggDg+fPn+P/snduOHMeVtdfeEZHHOveBoqzBLwgeX9DA3HgwN3Nhv4SeZ6jn4UtoHkCYC2MEjGEMNIBs2aYlkiK7uyojYu//IiKrs1uURMmSOknFB6Sqq7qpzjp0ZmSsWGsBwIcffkh/+tOfCAB+85vfAACurq7wb//2b/j444+PR6L/+7//o3/+538GADx79ozeffddvPvuu/j0009ps9ngnXfeubH7APDXv/71+O/v3bt3/OZUrDk7O8Pf//73G0e809NTfPHFF8fHnj59Stvt9vi7R7EFADabDZ49e/a1R8z1ev3NL9Ar8uzZs2/93mq10qdPn2K9Xt9wjHzxxReoqgqbzUYB4Je//KUCwOPHjwEAZ2dn+te//hX37t1TAPrpp5/inXfe0U8++QQA8O67704/C/rRRx8BAKbCRu6Q0XzymMUB6CeEHjx4QB9//DH/3//9X9X3fdO2beu9X4rISkS21tqdtfa07/uz3W53sl6v11VVtWbMSisU7pij6yPf8ng/OzlSD4gH9gfo4QDNtzgcwMMBOOxhctl5FQKM3n25KiG5QMwwQKLAi+RVrwQlToWwbKGci9FdBVNXyQVSOVC0IGNAoiDOE9OvgfNjynXXB03msF6nZ/DzofSyFAqF74IC6Zw0EeeVGWIdogKRGCwKzSII7ffA1RWkXyD6kCZ+okBjhIqk+EvVFAupCkYaCxQKPyYEwKjCqaY4UmNgqiqJH20H6jqg6yBNi1g5eGvhiRCY4VURVNPnPUdgFQqFwpSvc4Dc3grzQVUlxhivrq4OT58+vXzy5MlFVVUXy+XyEsChqiofQoh938fVajWbQ38RQArT8u4blqRRGPnP//zP49X+KICMPHjwAACOoskvf/lLAMCnn35Kn3zyCd59993bwsfx1wLA559//lIB5Ozs7MYPP3369Phz4+/Y7XYAgE8++YSY+SgyWGvpxYsXAHD83ZeXly+dsbh///7LHv5ejK6Nl+Gcw5///Gcws1prsd1uj+IFkASPP/7xj3j69CkA4PT0VIGbr0MWPwAA77zzjgLAu+++Oz6k09tb75O+//77N0raf248fPiQnjx5wvfv37feexdCaKy1fQhhCWAdY9zUdb3bbDYnb7/99snJyclus9ms1+t1U1VVEUAKs4Gyq4EUgOhRFCERUBRoTGXhFGMSREKA+FSwSnkSJfWH6DxWjE5X1auCshsl7X+Eeg/1HuQD1HsgeOiQHoMPgAs5DksAYZBJ4sdRCJnDc3wFxpjFaRF6mWefB1/nArn9MyJSxJFCofAV9HY/Ve5DYGtTObQoKESQD0B/gA4D4n6PSAy4CnI4QIYBGtL5nWOEkQgnEU4EXATzwo9IWqiicDFChwESAkQ0dbjlCKwUfdVAKodgTBI/iJL4AUVEWdZRKBS+nq+LvirCx7whIgEQmdkT0cDMA1L/x5A7quNYgP7RRx99ZS75LigCSOFrmQoj42PfkNmWbAX5APW73/3uW//3wLWA8m388pe/PIos//Vf/3V0pwDXIsCHH354nHm4/ft/SKHj6/i23zF+/8MPP8Qf//hHAMDvfvc7BYBHjx4dfy47Nb6Nl/7Mz1nk+AbowYMHdHFxYZ4/f26JqK6qqg0hLFV1ba3dichJ3/cnowCy2+22q9Vq2TSNtdYWAaQwCwjpGMspBHE86II0iQcaI5BLVJEnShCSmEBRkkiiWfiY5ZEiGdlINO1zFnDUB2hI8V46eFBMwgiFAA0RcJJeAxpjqsdy6nnHE01jsFIUJSF3/+XH7nDnCkemq9Km98fHysVZoVD4NnSyCRHEGCgbRElODgkhCf3DAMlRlsoMcRXC5SXk6gqyPwAhgGOACx4IKSaSRXAjPbEcjwqvynhe+5rHr78mGChqEYgqxDCkcimuralBTQ2tK0TnEK1NhelAir/SVHouKvMcehYKhTvnZX0fInLcyjh7fhCREpEyczTGBGb2zDw45w7OuSFHYMUQgg7DoL/61a90DgvFigBS+KHILu9X/lD/1Eexl+7YD3kwnfFz/zlD77//Pv/lL3+xV1dXrm3bWlVb7/0ixriuqmpX1/XZZrM53263Z2dnZye73W692Wz6vu8bytz1kygUgCx+JBnkWISevwGNkgrRQypFxyiGSMxF6SHFZMlXdO15MbpZRI4CjgQPDD6VtIeAOAzguk5CT0zPL0WBIXWBKKCUXieMgs+M/4yngk1hnrxM5BjFjzmLbIVCYV4oERQKJUJQgNiA1OZYxwFoG1DooSFksYQRiBHSKQ4YGOyz01FH94fCSIrCKnFYhe+KIBeUUxLnMEY9plxRgBlkGODUucZdC+paaNNA2wZoakjdIDiL6Cw8AR6KACAqEEQgyOOycq4sFArfgqoixnij/2N8vDAvRgGEiIIxZjDGHAAcmHmw1voYY6zrWuq6/tqu5J+aIoAUfi58nWPip96Pwk8Hvf/++/zrX//aGGOcMaYWkXYYhmWMcQvgrGmat3a73S9OTk7+abfb3dtsNqer1WrRNE1duj++mTLpdxdkp8D0kdENooCKZrEjb3IthpAooDKf6KuXkZ0sUzeLji6QGKA5zgveg4KHDgGoAiAClRTrpaogZgCTCesZH+ev3R9jBBYfeybK+enumbo/pu/J9PhXjoOFQuFVOAqmRIia5pdHEQTOgpo6OzYD4H06tykgMaYOEFUQG0QabfcCpbQWwAGoRG4ujigUvoVUTk4YiOCZEZkBk4QOGAt2FmQt2Dmwq2CqCrpZQ3cnkNUK2nWQpoY4i2gtvGFEpOLzoLn0HHkRAWa79KZQKMyAafH5eH/qACnXRbNDVVWJKGb3x4GZD865PREdAPi+74Oqymaz0dxZfOcUAaRQKLyRPHz4kH7729/S48ePzd///nfHzDWANoSwjDFuROSUiO4tl8u37t+//9Z2uz1bLBabuq5rY0w5NhZmCREds8STYHAtghw3EZDKdZeGCDgXptIYnTVDCGOcl4BFUtRV3hBuCiAYArhOvSbIkz6McXXt9YS16owFH9zcz+uBPR3juwrz4LYDZPp+FTG4UCi8EkQQJKEfWQQ5Zjcyg6yFVg6macAhQEUgPgDDkArSJUUIERRRFUASQBQEBMCqwpRjUeHbmPZaIXV1DGxwYIa3FsiCB5wDufR5tE0DbhrYtgWt19DNBrJYQNsW0VUQZ+GNgWfOhefXgsd0KxQKhW9iFDtEBDFGxBhvPF6YF0QkzByttZ6ZB2Y+ENEohPhhGKKISAhhNqeCMslXKBTeRAgAf/LJJ3YYhupwODTGmG6/3y9VdRVj3MQYd0S0M8bs2rbddF236vu+IyImopIi8BJeloFf+AnJqU6jgjEmN19HYWUxRATsB9BwAA2pUNWEgCpGmJw3PsepdQLAqnBRUHGEcISPASIRKjEXvAcgShJDQgSFmMrgRZNogHGj5Ai54+f0bYx/S8z8FYdBYV6MF2RTMaSIH4VC4VXRSRxjire6/h4zp9X2sUrOj3x+Ux/AWfynGAECNBWCIaZ1EGAFrAhUBKpxluf3wrwQpLirQARPBgMzDsbCWweuqlRwXtfgtgHaFmg72L5D7DrwagVdLqF9j1hXiM4iGIZPOhziuI0FxuMvnXkcaaFQuFum4sfU+TF1hBTmw7QDBEAgIg/gAOBgjBkAeGttrOtahmGYzZtXBJBCofCmQQ8fPqTdbmdExDFzY4zpvPcLAMsY4zqEsI0x7rz32xjjkog6Y0xljHF3vfNzpUzIzgTKq8+nEymjs0MVLAITI+zhAHfYg68ugRBAwcMGj0rGzPD5QQpYCBqJ0JhypyEGh+z+OMZixZj7TOS6+2TSizK6ZIjo6A6Z5zNO3HYXlGLt+fF1DpBiyS8UCq/MeM7OThAASaZnSt0K1oJcBGkF+ADKIoh4D/Y+TQJNzvuqColZ+Ih8LKue9xmvcNck7xDgs/Nj3IJNMVbqHLiqQW0LbVto34H6BdB34OUSuuihfXZ/VFUqPTcGgQgBt6Kvxq2IH4VC4RWYxmCNX5drolkzlqB7Zh4ADMw8qOrQtq1X1bjdbuXPf/7zbN7AIoAUCoU3ihx9xX/4wx+Mtbby3jci0qvqEsAawEZEtiGErfd+FULoQwiVqpbOj1egDEBmRHZy5M5KgAADhQ0e7WGP5vIC9vJFEghyDJYVgcE8HSAMhVOAYgATwEQQa1KBZo72gmp2g4zxXjF1hhw/l9fih6qkW2D2MVjT29tfF+6W6TFvmkNcCtALhcL3RVVTHFZ2/olhRCjIubTAoanA2flIwQMxwmTXB3B9PiSJUBGA/XWcVjkkFb4BARCZMbDB3hgMxh4FEM0CiNYVtE4iCHc9qO9AfQ/qe6DvoV0LrWtoVSEYA0+EyIyAa3fJcdU2UMSPQqHwjdwuO59u47GkXBvNi9EBQkSRiAIAb4wZRGSw1g7DMARVlRij/uY3v5nNyKQIIIVC4Y1AVQkAffjhhwzAxhjrGGM3DMNaRLbe+52InDjnzuq6PrXWnpyenm6Wy2VfVZXjsYW4UHgdyMoH8aScOU9+MBOIUicGQ3P/R4TJReFzHT6mHg+FU4WKIIrAiIAkOT9SqXvILpAASMydJ6k7BGMxbBZBOK+yneME9VT0uB19Nb5/058r3D1TC/5t50eJBywUCt+JLM6PqZZCQGAGDAPOAlIngUP12N+VVwZAiEAiqRcEBKcCM/OOr8KMoPQZCmzgjcWQHRxiHaiugboGdx2460BdB14sQIse1C+gywW07yFNg1BVCM4hMB/dHzJuE/GjOCULhcKrMhU9pr0fxQUyP/KxXZj5WIIO4EBEB1UdFouFDyHE/X6fohpmsjyjTPgVCoXXHlWlR48e8UcffWQA2D/96U9V27a1974PIaxFZAvgRETO6ro+3e12J2+//fbu/v37q5OTk65tW2etLaPzwmvBcdKcb44kjoXahiGuQqgqSFUBzEcxhKZl6XNjMtljVGAmxe2j8wOSb1UgEo/xV7fHVGPq9NxL0KckDeumMFK4W24LG7dvR8pFWaFQ+L4oUepMIEIwJkUKVQ6hqqBtC3QpeoiXS5jlEqbrYJsGzjAqiahigIvx+vxeKHwDacREEGZEYxGNS+JHVQFVBWqa7PzoYBcL8GIBXixByyWk7xHbFqGukwBiDYJJAkgEjo7dafRVGcsUCoVX5Xb01SiEAGWsPTeISJEisIIxxhtjBiIamPlQ1/VQ13VYrVZxGAZ99OjRXe/ukeIAKRQKrz2PHj3ijz/+2AAwdV1bZq6MMW0IYYkUeXWqqucxxvOmae6dnJyc/eIXv9ienJysVqtV2/e9tdYWQbjw+pInz8laqKvg2w46DIgS0YLAmtwUrxPJrTLZsghCueyVcgQIjhfYWQCasctlyihyjAXozASRcYL9jneucOT26jMRgTGmFKEXCoUfhDyDAFEFkYFHOt64BlBjcj+IAVkDZQJLBO+v4AhwEmH8ABs9jMprce4r3DUEJYKygRoL2Ly5CqhqcNvCdB1MFj9opEi0AAAgAElEQVTMcgFaJOeH9j1iUyPYVHw+uj8iUvdHLOJHoVD4B5iOqW93gRTmhzFGcgSWBzAYYw7GmKHv+6FpGn96ehrv378vDx48mM0bWASQQqHw2jI6P/7yl7/Y9957z3rvqxBCdXFx0Q3DsD4cDltVPbHWnlZVdbZer89PT09Pz87OtmdnZ8v1et12XVc554iIigBSmD2qevQ6XNdeEIgYnOMx1BhE5wBXgV2DaA7Q1/XjPQocItfl56pAlGs3iMgx+oN0DBSh10BF0Bx1pem9wzQSKz0+E7fwzxZVBTOjqir0fY9hGI7ix9e5QQqFQuG7IkDuSVDAMBQWEQATwxCBx0UOouAQwZdXMG0HbmrwocrnRv8anPcKdw4hiWrOgqsKXNeAc8foK9P14K6HyZ0f2nVA10HbBjI6P5jhOcdeESHm4nMAybFbxI9CofCK3O78YGY452CtRd/3WK1WqOsa1pap6zmR+z/EGBOstd4YM6iqV1VfVVU4PT2NuE5G1OwYuXPKp6hQKLyWqCp98MEHZrfbmaurq2q9XleXl5etqnaquhiGYee9PyOi87Ztz1er1b31ev3W2dnZ2cnJyXaz2XR939dVVZXjYOH1YLygPE5wXK9AJ+DYC6LMUGsAaxGtgTBDX8cL0bSEMDs/ksgxFrofhRFN7hDItROEJkXopCleZI6TQrc7JJIGGyeP0xx3+2cFER3Fj5OTEzAzXrx4gaurK3jvj7b82/+miCKFQuFVGY8WowhCRIgKwFowK8J4jgeBYgS8B5ZL0P4KNBxyPwgDlxdQ7/NCgELh5aQIVQZZB65rmLZN8Vd1A+57mOUSvFgAx8LzDtq2kLpBrBy8MfC58DxAcZzhmizQKeJHoVB4FaZi6SiAGGNQVRW6rsN6vcbJyQnW63URQGZGvtZRIorGGJ97QDyAcDgcAoCIfDU/F/EDKAJIoVB4PaFHjx7xbrczxhi32WzqFy9etDHGJTMvVXWjqichhHMiOquq6uzk5OTs7bffPj85OdkuFotF0zS1Mcbc9RMpFF6V2xeUt8uzr7+RhZFRIPlpdu9HYIy+EkCz8CEKjTn+SgQqExEkw5RFj5lHfo1zVDcnzG++n2US4W4Z3R+r1QrOOTRNgy+++AKff/45RAQhhK//OywUCoXvQhbrRRUxT1JHCNjZY78HhRomdBA/IMSQooyshTUGFDwohLt+FoW5QwSwATkH0zSQrgdXVer9WCzA/QK8yO6PtoE2DcQ5iLU3Iq+S8EGIIhCd93irUCjME2b+iggyLjy6f/8+Tk9Psd1ujy6QwnzIDhA1xkQiCjkGKwAI3nv5+OOP9cGDB7M7ORQBpFAovFZMY6+urq6qzWZTX11ddcy8UNVNjHEjIifMfLpYLM7ruj7fbrdn2+325OTkZLNerxdN0zTGGMNj7kyh8JqhOR1pTFu+7r1IcVEcA2zwsNGDR/fE68TU5CIKkuzyGB0gRyfIdfyV6nX3x3QF/rxX4yeXx/UE+vXjZTL97iEiWGvRti2cc4gx4nA44OnTpwC+PuO8uEAKhcJ3YozUA5A6GhRChKAp0lGNAVxasY8QQYsFoqQzPwFpUcDhABADfkjrIMaIyHEMUI5JP1+IUhSqYUhVA22T4q5yr4fWNbjvga4DL7Lzo22BtoXWNaJzCMbc7PtAzjVBCessFArfnduLh8axMzOjrmtst1ucnJxgu90eI7EKd4smJMYo3vvhcDgchmEYRMQDCKoajDHxcDjIv/zLv8xO/ACKAFIoFF4jRvHj448/NmdnZ26z2dQhhJaZFzHGdQhhq6onxpjTuq7P+76/t1qt7p2enp7udrvtcrlcdF3XOufcXT+XQuEfRZMCMrmX3BIsAus93DDAHvYwIYBn7oZ4KVn8wBh9pXkiZ3R/TDtBNHkn5BgLdv3/yKnqs2I6Of7VKCygTCnMB2MMjDGo6xqHwwFN02A0D75MACnZ54VC4TtDBFEFE6UKKzAECjIMARCQjjnGOaCp07kPlP4dCBIj2HtE50DDAA0B5APID2A/ADG+fgshCj8YSgw1BlLVkLaF9D3Q9Snyqu9BXQe0be78aI8CiNQNonMQ51LpOVGOvSIIkLo/MOnDKue+QqHwitweL4/XRkQE5xy6rsNyucRisbirXSzcQlUlhBCz7nF5dXV1sd/v9zHGgZl97gOJu93uqI/PKf4KKAJIoVB4DVBVAoBHjx4xAHN2dlZZaxvvfT8Mw4KINt77bQjhTETOqqo6b5rm/Pz8/K1f/OIXb223281isVi0bVsbY17TNui74/bKjMIdkufFx/Hi9W1aBZrEjwHV5QXqF89RXVzADANY4l3t8fckR1uNIogoKN4WPrL7Y1zZqsCYlD51g8yV678lncQojV0ghTky5hPHGCEiEBHEGGGMOR4fp8fJIoYUCoVXhSiFORJRdncAYIYCMDZL4lUFUoCVwLnxSoggDARnQRcX0Ks99DCAry5hLl+Anj8H6WH2sZCFH5Hs/AirFeJiibhcAv0SZrUEd2PcVZv7PhpILjyPY+m5YYRceh6R+j7i6EHO58UifhQKhVfhduTVOG5W1ePYeuzYK/MO8yLGKIfDYXj27NnzZ8+ePb28vHwSQngRQtgbYwIRRe+9/P73v5d33nlnloOOIoAUCoVZ8/DhQ3706BGdnZ0RAH78+HG1WCzq/X7fxRiXxpjV4XDYquqJtfasqqrztm3vbTab89PT09OTk5PdcrlcNE3TWGtL7NX3pEzizYwbBoHraAuS7AAZBlTDAW6/B2XnxGvJWHR+FDnSpiLXsVjZ5QG6uXroWIo+KeacEy8TFMe/M2bG69ze8qYyvmcicj3pg69eoBWxuFAofC/y+YoomyCRy6WJYIwBWwWrIubzIicTCIQJMAZoO+BqD7m6Al44gAkcBSACYz9xTZbj0xvBOIkIQMbFSsC124cZoCR+SNdBlivoag0sl+B+Ac2xV9onBwi6DtrUkKqCVNUx+ioaRlBBgOY1KYpxVFnEj0Kh8KpMxY/pWPn24qHpWLswH7IDJFxeXl59+eWXF19++eUFEV0R0TAKIMMwyPn5uQCpJ+Su9/k2RQApFAqzJUde0Xvvvce///3vjTHGnJ2dVVdXVw0z9yKyFpFtCOGEmc/quj5frVb31uv1vZOTk9P1er1bLpervu9bW4IjC28iUyFkLEkVgQkBxg8wwd/l3v0waBJ2NEdh0RiJNU5Ci0BVrid0VHHs0Ji98HPt/piWaU97QQrzYXpRFkI4uj9uCG/AV+4XCoXCKzFOAuVjRxzdjFkVIcMg2OQCycIHcXpcjQHXDejqCnpxATEmOURiPg+qgvwAKnFYbxQCQIgR8/ouUoVBPv8YA3EVtOsR+wV0uQJWK/BqnSKvFgug6xDbBtK2yf2RI6+is4g2iR9eFTHHtEn+nUAefpbzXKFQ+A58XQwwgK8sMCrj6HmhqhpjDMMwHC4vL6+eP39+6Zw71HXtAcQskMgf/vAH/Ou//ussBxplQrBQKMwV/uCDD/jBgwf8v//7v2a329nD4eCurq7ai4uLhYhsVHUXQjgNIZxVVXXW9/29e/fuvXV+fn6+2+02q9VqUde1K66Pws8KnaoirzEpW+GmsHEsP9drdwgAyoKBAEchQbMQkhvS7+xpfB1Eyekx2rzH/g9mRjlkzZPb7o8xAouIwMwvXclWKBQK34lbIggASD6PMTMCFHAGgMsnkhSd6JhB1gLGwHCKUlQAkQhqLZQZ5uIF6FDisN4khAjeMAaTpnWMCqoQwMYAdYPYLyGLBXS5BlZr8HIFjL0fiwW0a8FdB6krSFMjGoPAfN35MRaeH023pfOjUCh8f142Rh7H1dNtfLwwH4ho7PSIzOyZ2RNRiDFGIhLnnNR1rb/61a9m+8YVAaRQKMwNevjwId2/f99cXFzY58+fW1V1quqqqqqHYehFZHU4HE5E5NwYc9Z13Xnf9+fb7fats7Oz83v37u1Wq9WyruvaWmuphOoX3nT01u1rDuXraqMKq4KQ82B1InyMgsgogkxFjuOAeY4N6BM0T2gx8y0XyMx3/GfMKHqEEG5kFZeupEKh8IOR+0CyHfAYGxKgUGaQTYI5GQZx2oxlsGEQG5Ax+SSaHQDOAbmrCMygQ564njhHj+fVwmuFMiMYi6GqADawImAeYKsKaDvE9Qa6XgPL7PzoO6BPBeja99CugTRNEkCqCsIEASGQIoAQKYsfuDYdF/GjUCh8H6Zj5elj0x6QIoDMlzwWESKKROQBeABhLD+31koIQR8/fjzbN64IIIVCYRaoKn3wwQf04MEDevLkCW+3WwugIqJKRGrnXL3f77sQwjLGuIkxnjLzmXPuvO/7e8vl8vz09PRsu91u1+v1qu/7zhhj7vp5vUmUQcjMeYPeHgLAUDhVVHmCOeTccxmL0UeHCJAvxLNooJomhKD57jxfmDR/wFB9mYOg2L7nyPj+xBiPIoi19sZn7GVxWOW9LBQK34tRCEGegM4TRZEURBbMks8fhGg4dYUwX09OGwO1DpQdIRBJQoi10NFRGQI4BHAMJRrrNUMBKDHUWERXA8aCgNTfUdWgxQKyXkNXa9BqDc3CB/VdLj1PsVexqhCrCsEaBEozWjEXnUcAEQqZTkiWc1qhUPgejGPi24uGbhejjy7rwrzI7g8logggEJE3xngAkYiiiMx+EFEEkEKhcOeoKgEYXR+mbVvz5Zdf1sMwNABaEWkPh0MvIkvv/TqEsBmG4bRt2/O2bc/feuute+fn56e73W632Wz6qqoclRmnws8IVcVYm/0mfPAJCieCBhGIDBMDrkLAQQQiEdPi96MTBPn5TwrQ58r1vmke/AOpt4TBbABQ6QGZIdPYq+l2u8fldhdIoVAo/ENM47AAxPyYEmVHSJr4tkpQJZASmChFYlkHGE5F6dZC+h7YX0FDAIYBdHUFt78C7a9SSXrhNYIAYsBacN1A6hpiLQIztK5BfQ9ab0CLBahfAH0HaVugbSFtdn04B28NAhM8ETzSYpOj80P1psm4jEsKhcI/yCh4TB3UU9GjdIDMkxyBJUQUiMirqgcQmDmIiIQQZO4iSBFACoXCXUIPHz6ksesDgHXO2Riju7y8bEWk9973IYSFqi5jjBsR2QDYOed2TdOcL5fLs7Ozs9N79+6drNfrdV3XzjlniwBS+NnxBn3ix/TyWiNIGCwRQQV+0v+BsfhcR+EDIFyLH8dL9iyIzJMk24wxWADAnFbzlkPY/BjFDWstrLVH18540TaaDovwUSgUfmhutHuN54ccn4iYziVRCRZILhCThBF2DnAWcBZS18BlDxz2iPsDcHUJdi6diXIMVjp8TRYYTHfgltWUbt3O91w7Y8bJP7zMyEvHF3eM+qTJv1NjoM6B6gbUtOC+B+oaYh3QVDD9ArRcgvoO1PWp5LxpoE0DbWr40fVhkgAyIJWdJ/HjuvBcJyJIoVAofF+m1zZT8WMqfBwjj1HG03NjGoHFzIGIfI7CCkQUrbVS17U+efLkrnf1aykCSKFQ+KkhAHj48CH99re/5cePH/Onn35qHj9+bDabjXv69Gk9DENjjOkALPf7/QrAWkQ2IrJj5m1VVbuu67a73e7k5OTkZLfbnaxWq/ViseiZuWgfhTeeGyWUU96gjz4DYFVAY5pcFgHl6CuN49c58opwXYgOHOcMiChN6NzpM/lmpjbwtHHe3qA38w3BWou2bbFerxFCOK5eA64v5KZxZiUGq1Ao/FAo0nnthkcjH2sEqQvCMkGYYAzDGgPjHLRyoKoC1RW47SCXl9D9HnJ1BVw0UOfA+SQpxkBFoDEez6+q1+faqfNyPOcykgN1dKEWvhuKa1eP5MgzxWQRxHheUQWrpHERMdTa1O/SdtCuBy+XkH4BZIEDbQN0HWjRg7sOaLL4UdeIziFUafPGIFB2f6giqkCJUuSoSOn8KBQKPxi3x8PTvo+p8FGYJ1MHiKp6Zh5UNQAI1togIhpCmPWbWASQQqHwU0IPHz4kAPzgwQN+/PixAWC2261VVXd5eVkbY1pjTBdjXIQQNgDWMcatqm5ijKdt2+4Wi8X23r1723v37m13u91qs9n0TdO4LH6UEXrh5wNlMeRN+9RPBsBJ1BgnXnJm+TgxEyMIk1L0HClFGH/kWiia26FhnDyf7luJUJo3VVVhs9kghICu6/D555/j2bNn2O/3R0HEGPOV97RQKBR+CEYRJIdwp0lzpB4IEKCUHldjAGMA56DOwVQDqHKAq8DOQaoK5BzUJKdIZIZUDuHqCuIDJHhojNAQoRLTeXeyUXaDWBVYVVR6HUNZ+G4ogABgIIZnRkwlYHlLBfdMBKOCKgQ4EZAxiE2DuFgidgtodnpw14PaFtw04LYBZwFER+GjqhCcQ3D26PzwRAgEBFUEZNfHKHyMO1nOY4VC4R/kZddkt8WPqQNkjtduP3fy+6VEFJjZAxiY2RtjgoiIc062263++7//+2wvYIsAUigUfiro/fff5/v37/Nnn31m9vu9aZrGhhCciFTMXMUYOwBdjHFBRCtr7Y6ItsaYnapuQwinTdNsF4vF9uzsbHN+fr7abrfdJPbqrp/jz4YyMXtHXFdH3IhFoJf9zJvCsez85ipUFUkPZUEkrUSlyepYne3n9GX7NT1+jQXb4zaNyCrcHVVVYblcwjmHpmnAzDgcDhiG4aUXbKOYNdfPYaFQeP1I0w8KyWI/pfzHVIdFDCGGGgWshcYAW6X4K1h7LECn/DUMQ4xBZE5iSXMFGYa0HQ6pJyRGIERI8OlrkRSXBcBJRK0CI5qcCYVXYxJ7FUEIRNizwcCc+juIUrxZ7ncxRHAqSQyJEeQcYr9AWG8Q+yW070FdlwrO6wbUNOC2TdFXix4yih/GIDibXB/M8Cb97iCCoAqh686P42Tl3b1KhULhDeV21weAGxGzxphy3TNDcgm6EFEc46+mEVjOOfnb3/6GBw8e3PWufi1FACkUCj8Wx2jg999/n37961/Tbrcz2+2WrbW2aRoHoFLVGkDjvW+z62Ohqitm3nRdd7JYLE4A7ABsvffbtm3Xm81mtd1ul6vVqu/7vi7Oj8LPDcJLhI+vfPcNQzU1cqrkFanxVg+IQrMbhCYTQ+Mge65MY5PGgu3D4YBnz57BWgsRQV3XqKrq2DFRuBvG3o+6riEiePHiBay1UNWjUDV18Uwv7MpKtkKh8EOhOSoJSNFTCkCZMDZEqALKCmcYGmMSRSjFYpHJ4kfuCYExgLWI1kFdhbjfJwHEOiB4yOCh3qe+CT8AUUCaRBAQwUjMMVmCMl3+aiQ/K0Fy9NRAjMEYDGzgmVOxuTGANWBrU6cLAOsCjArYVZDlCnG1hi6WQJ+dH20LalqgrlPkVddC2xZSVYiVy6IHwxOn0nMoggoiFBGKnDJaRPtCofCjMB0bTyOviAhVVcE5h77vsVqtUNd1ue6ZGUSkzCxj/weAIcYYnHOxrut4cXGhp6ensz6BFAGkUCj8kIwRV3jw4AF9/PHH9Oc//5nquubVasV931vvvRWR6urqqgbQHA6HLsbYA1iEENbe+1UIYbVer3fb7fb83r17Z23bbo0xa+9975xrm6ZpN5tN03Wds9aWM+OPTLkQek140ydXVaGaV9nnGA49xnFkcSRHQ4zZ5KMzZI6vzHQyfPq19x5Pnz5FjBGXl5fY7XY4Ozs7xisV7o7xPTDG3ChBjzEixngjy3j8+SJ6FAqFH5MxqmjsaQj5PpggkgrRrbMQIohhEBPYMGAIsGmSfRqZRVUN2l+BrIUOA9QcoMZAvE+CSUgLEFQEEgI0KlQIOmZzFb4VBSHkyKuBDQ7M2ZVhIMcCewdyFnAOMCY5dQAEw+CqBhZL0GoN6vvU9ZFdH1rX0LqG1FWOvqpS54c1GCg5PiIDXgUBSK4PXJeeFwqFwo/FNAZrGnk1OquXyyXW6zV2ux1WqxWcc3e8x4Up+T1TAJGZ/bgBCPv9Xpxz4r3XDz744K539WspAkihUPhHOLo8Hj58eBQ9APBf/vIXWq1WfP/+fXr69KkhIkNE7ssvv6zquq4Ph0M7ET5WqrqKMW4BrIloXVXV6XK5PD89Pb23Xq83VVUtVNUSkWVm27atcc4Vb+RPRBFB5sxkiv9YmplWiILGtaGZ1/J91JsD5TGCQ0c3iBydIKPoMb4e1/fnxbgCarxV1eNk+jAM8N7j+fPnOBwOiDGi73s0TXPXu124xejYGbfbq9kKhULhx2Z6hhNcnwJVU7G2IUodH44QmWBypCIzgZgBJhAbEBvAWHB2iCgnF4IxBuIccDhAvYH6FIVFkiKZdMiLEqBjPlfesfmde+eCEhCZcGCTnR+pkwPWpvfBpugrWAeMJfZVBbEOwTlwXad+j34BtC2oS64PbVqgqaHOQeoKMYsf0Vp4Jnikz0RQSQ6ULHqMsVeFQqHwYzGOi6fxV6MAYozBYrHAW2+9hZOTE2w2G7RtWwSQeaCj8CEioqoRgBeRICKemUOMMaqq5IisWVMEkEKh8F0hVcUHH3xADx48oCdPnvBnn31G/+///T9+8uQJn52dcYyRrbVmGAZzdXVlAJj9fl+JSEVE9dXVVRtj7FR1AWBJRCtVXTvndk3TbOq63ux2u912uz1brVany+Vy0TRNp6o51YaImYmZywxToXAklWYqG4irEF0N7w7gGMGaBYPXkBt7nZ0eKqkAXWNMueM5f1xEb8SD0VgkOtPnfnuyfHQTjN0fzjksl0t47xFjvMtdLdxivGgb369RBLHWHr8/RmJNxa5CoVD4MdA8mT3K/0IAE43mSCgRLBGUGUwpOosBMDGUTeqbyE4QchZsDVDXkMMBNBzAlUuOEO9BMYJiBA9D+rlDEkY0eFAM131dhW+H0utuqgo6uj6MAWfRg52DaRqYugKqFG2VIq7a9HXTQJsaVNeQuobWo1BiEaxFtAaBgcCEoIqoighAoBCk8VQJLysUCj82t10f02seAMdrnvV6jdVqVXpAZoKIaAhBDodDPBwOh4uLi8Pl5eUQQhhU1TOzt9aGqqoiM8swDLM+nRQBpFAovCr08OFD+u///m/64IMPCAAvFgt68uSJ+ad/+icDwDRNY4ZhsCEEC8A555yIWFWtYoz1xcVFLSItEbWq2gNYENFSRFZEtFqv19vFYrE9OTnZnp2drU9PTzd93y/qum6dc9XdPv0CUHLs544SIxoLX+eL4uBhDgdY72H09Z5A10kB+rilKjZNK1E193+IgswoeuQx2Iw/s9POCGY+Ch23XQXl725+jN0fIoIQwo2Lu/H7RfgoFAo/CeOxhggxOyKVKE1uM6XTZr5vrIVRBROBOZ17iBkwqTCdqgq2rqGHA/hwAIYD4D10vwdCAIUA9QEueJhhAKoDdDgg7q/AhwM4+Dt+MWaOAqwKl92rbBihqiB1EjfIOcA5cF2B6jo5PpoG3LTgJn0NVwFNDdQVtEpOD3EOWlUIhhGtRbQWgRmRc9m5KiR/PlIPyXWEWqFQKPxYTK9jxnHy1EEdYwQRwTmHqqpQVWXaZy7EGGW/34enT5/unz9/fnlxcXGx3++v9vv9HsCgqt57H6qqCsMwCAD9j//4D3348OFd7/pLKQJIoVD4No7CBwDabre02+24rmvz2WefmcViYQ+Hg22axomIE5FKVaurq6sGQL3f76sQQhNjbESkFZFORDoAHREtRGShqgtVXa3X681yudy8/fbbu9PT08Vms+mapqmMMeVYVSh8I3lQyQbRWgxNC+kXEBE0AFgERl5vAeSG+CECjbn/I28s6XsyCiH5n9FMHSDTC4FR/FDVFDeS83DH1U9F/Jgf01Vso1A12vpvv19FBCkUCj8JExEESNFGx6MRU0qpYk6xR0gOEMMENhZsGFw50FCBmgFmGKCHATQMoOEADAPocAB5DwweCCE5QAYPCh7x8gJkDDT3c1FxLX4tDIUTAavCWoNIgK9qSN9Duy4JIHV2gDRtEkHaFjS6P6r0fXEuxV3lmCuxBtEwojGIxiAQEIBr1wddx14dBfs7fi0KhcKbz23xYyqCjK73cSxdmBfee728vPSfffbZ5RdffPH82bNnz5n5wlq7t9YOIuKdc56ZY13X8j//8z93vcvfSJlULBQKIzku/zre6uOPP6b79+/TZ599Rr/+9a/5/v373LatiTEe3R6Xl5fOGFO9ePGiHoWOGGMTQmhVtQHQMnNb13Xf9/2ibduemXtVbUMInYi0McZORLrT09PVycnJcrvdrlerVdt1XcXMTETF/1go3IBu3Y53KRVoOgdUNcjViGYP+zpPoKd21zRxI6kDhLL4oTECMYJFAIlAFJBRgBRj+tXYDTLXi/zp5PgohBhjjo8dDgc8ffr0KIzUdX0URwp3hzEGTdNgvV7Dew/nHKy1x/elFKAXCoU7YZxoynf11mNCqQdkFEAiMywbsDEwIcBUNagJ0GEAe38UOdgPoP0B7D3Ie+jgQcMA+AHkPaiu09gDAOwVdH8FCj7lb42TWtmBIkRQoq+6D26dqOllD37Dz3/jy5L/wRj9Ne0IG/dFJl+/6v/x+ssxfCxFcvIoRHEumR9dNjmudFzcQFUF2y/A6xV0sYR0HaiuU+9HXQF1k4SPtoFW144PcTZto8vDGERmRCJEQr7NGxRRJD236QTkq798hUKh8L247WIfFw8xM+q6Po6ll8slqqoqY+eZoaoyDEN88eLF4cmTJ/unT59eNk1z1XXdvqqqPRENAMIwDBGA3Lt3b9anliKAFAoFqCqNoseHH354o8T8yy+/5LZtebPZ8MXFhTk7OzPee7vf7x0Ax8xVCKEWkRZAC6BT1TbG2McYO+99Z4zpu65bnp6erne73aqu6x5AE2OsY4xVjLEOIdTL5bI7OTlpl8tl1zRNZccw9UKh8BK+KoKMEx2SC03FGCjxrCOgXomjCDJ2gEgSQaKAVFIha0wukDSozuqHKGn4+GkAACAASURBVIjp+t/O9HUYB/vjpPk4iS4iuLi4wN/+9rdjOfput0Pf90UAuWOcc1gsFjg/P4dzDl9++eWxtH5KcX8UCoW7QpGPQUCOPaLjJD8zgWFgmAGTSmjJOVAloBhAoQYNHhw8zJDcHqYZwEMWPHwAhiH1ggwD4CpwnujX6gXIGujlRRJJxtJbJPHDM6dJe6JJd7pe7zT01vKO2/fTz32XUzohxU4ZKJzqtQiSf2UAEIghlPbxuCuTn7n5f8u3WfwgouPvsCpwmkriYStIXYOqOpecM0AMNgwwg+sa0rTAagNd9EDXAVWKvkJVgZoWWlfQtoZWNaSqoFn4EGtStwflDYAQIyBHXQEQleui8zwOKrFXhULhp2Lq/pjeGmNQ1zX6vsd2u8V2u0XbtijTP7NDVVVCCMF7P+z3+wMzH6qqOqjqgYgGa603xsTD4aAvXryY9emlfLoKhZ85Y7H4b3/7W378+DF/8sknfP/+fd5ut/zkyRNjjDGXl5cmhGCstZaIbFVVzntfMXOlqrWqtqraxxi7GGPvve9FZJFve2vtommazdnZ2ckvfvGL7WKx6Jm5EhEzbqpqrLWurmvX972z1hbXR6HwfZj1sOMfIIsfYwTWGH+FKKn3IwpUIkgNoAxGmoxQ0bER/a6fwdcyFmaPK6JGvPd49uwZnj9/jidPnuBwOMAYA+cc6rq+wz0uVFWF3W4H5xy22y2++OILPH78GBcXF9jv90cxa9oDUrpcCoXCT81UgI24dkQyEdjkSCTDUIvcraVHlyXlvg/2AXwYYLP4wd6DfQAOB8gYlVXVUJccC2haoKqOTk3KJbeaHQkHY3EwBj5HP6YZ+ewSGRc8AKnnKw9qpkfO0aMx/f74na87whIAo4paBUYjphcZgiR+7JkR8j5O/8+KiStk4vZI44q04IIolctbUdQSwDHAGAutG+hyBW07cN0kkSmLTciOXVPXoK7PheYNqKpSF0iTi82bClJXkKoCnINaC8lRVwGaxBsogqbbKEhCjipkoiull7lEzBQKhZ+e6YIgEUHbtthsNnjrrbew3W6x2WzQ9z3c6CQszAYiUiISZo7GGM/MAzMfiGgQEX84HMJyuYyXl5fy3nvv6ZyvdYoAUij8TFFVevToEX/44Yd0dXVlYoymrmvjvbfDMJiLiwvLzNYYY6uqcsMwOADuxYsXjpkrAPUwDE3btm1VVd1isVhaaxeq2nvvO+99PwxDF0JorbWL09PT9Xa73a1Wq81isWittXYUX0SEARARMTOztZaZeb5Hzp8Jt1dqFObOm/wnc7P8XHPpOWJ2f4TRASIQydETUQBOkyFZCnkttKExBouIEELA4XDA4XCAiKDvewzD8BWXQeGnx1qLpmlgjDlGlj1//hypE/Ca4gApFAp3zXgEGkcJx/LrHEWVvpdvFSCr8FGg1gDBAibAWovoHEwI0OABH4GmBh+yC2R/AGWnAioHWAP1PjlC3FXKewchECNYg4EYnrM4LNmdkMUQwnib914x8VxMBBH9qjgyvXdbNHEisBKzG0KuHSA5PjRYm9wpOXlXp9t0QmeMyaKJ+MEGTASFwsYIUUkiR9cD6y3Q9aA29Xuwc4C1QBZC1Dlw00Cr1PuBqkquj7Hno64Q6+q62NwyPDM8CIGACGCQmKKuNIkfo9vmRtzVjJ2whULhzeNl5efjNjpAVqsVNpsNVqsVnHM3FoIV7h4iUmYWY0w0xnhjjCeiQVUHa+3BWjsws7fWxqZp5Pnz57O+6CkCSKHwM2MUHQDwYrEwL168MMYY+8UXXzgRcarqXJLeKwBVLjWviage465yoXkjIq2q9m3bLs7OzraLxWJhjFkMw9B475sx2oqZ28Vi0W+32/VisVi0bVubkt/yWjBdxVyYM3TUCN68S1s9zkCoZMFDFRoDIEn4IIlgiVBR8FiMzskDwrn088jMXqCp0DheJIyD/7EYcL/fw1qLy8tLeO9LSeAMGLOL67qGquJwOKCqqhQjcyvSrBw/C4XCHJhGHzFRniDPj41uDE6T+4YZIpw6QoyBxBS7ZGKEjQINIUVhNR4YBqAZgKEBDV1yLVRpFa+0LfTqEhIjggi8AAOP3RSTaCaRowAyOlGO/VgToWMURY6nctVbQsdXT/Lp3yk4RojPvSTx+tVQYogxiNYh5E6NaYfKUSw6/g/z0oocZwXOAginY76HwhEBVQ3uF6D1BtRnAaSqQK4COZecN8aCKgetHNS65PBwFuIcxFnEvEnljl0fngmBGR7J1RNyyXnMBedHgWvyGl7vd6FQKPw0fJ0TYLzmcc6hbVt0XYe2bX/ivSu8KkSk1trgnPPGmEMuQN8DOIQQhuVy6Y0x4Ve/+lV89913Z52yWASQQuFnQhY+AIA/+ugjfv78uWnb1gKwT548qaqqqomoCiHUqtrEGFtVbYdhaIioUdUuhNCM34sxdiGEru/7ZV3Xq5OTk7PNZrPquq4LIVhVtSJiYoxWVV1VVa5t29o554q74/VjzlbGQkKPkwCE6TTBm8PE/XEj+iqCo4BiBGIAi80537ngFZPP70xLP6cT5tNCdGPMdVHq5G+w/D3Oi+n7N97eFj/Ke1YoFObEdGJcQAiqKTIJqQ/D5MJwywwDgiWCZYYVgY0CKw4mVuCQ+kG4DcBhSJ0flQPqGtFayHKJcHUJ9UnQ994n0UMiEON1SfoYcTk6PYEb3SE0OX9TdnROXSDjd77hCQPBp/9b8DhmgQFJGDA2xXY5l0rLcVMwOv7cNP6KU+cJmJObwyRXh1qL4ByoqYG2A/cLcNuB2hZc18kZkqOwkLs8xFmIsVBnU6F5vg2GEZkghhHy+xQUiDGmzg9oEj7y6yMi16JNEd8LhcJMmMbBAjcF2jJGni8TB0gwxnjn3GCMOYjIAcCBmQciCm3bxsvLy1F/ny1FACkUfgaMcVfvv/8+/fGPfzSff/65ZWbrva+urq5qZq5VtfHet6rahBC6EEI3lpiLSGut7eu67qqq6o0xrYj0IYR2tVot1uv1qu/708Visej7vo0xMhHReKuqzMxsjDG526Oc5V5Dbk/CFubL9UXvGySEaI7mGOOtRNPkSRQgRHCM0CjXLhDDINXrVa6ja2KmERDTvojx/jQOa/y6MD+mPR/j/enjL/uZQqFQuEvGSCQFJUFBFZp7IxjJncEAIhEMp44MywSnBtGmbgkTYxJArIEJAewcaKiODoZoGLHrEC6vIH5AHAaI98k9EgNMCKm/S1NXCFShMZ2raRRD8n7edn/Q5PERmvz35lcAiYBjAFkLIYKEcOwdUWuhVQ1qO7BzKdZw8jrdjsHSsfeDTRIxmFOvh7Ug66BVBW1aaNukAvSmTfebGlrX0CyAqDGIxqQ+D2shxiQnimEEc11wHjk5PSIlcSpKdnqMPR/j/o3ix6TwvFAoFO6S29c242PT8XAZG8+XUQCx1gZr7WCtPTDzYK0dYoyemQMRhdVqFf/617/O/o0sAkih8IYzih/vvfcef/LJJ+bTTz+1qloNw1BdXFy01trm8vKyI6LWe99l8aOPMS5GESTG2Flrl03TLDabzdI511trW+9907Ztt16vF33fb5qm6aqqau76ORcKhTdsMDmJxcAogowukBDAuQcE2QlCYsA68cLoZNB9l8/jJbzM2TEVPm47QIoIOU++7e+NiEp0WaFQmBVJBJHkYECKUCIiCPR4DpVcCm6OMUuAVYVkl6IxBsYaSIxgmwQGWAOxycEgTQNpO8gwQIYDdPAgP4C9B4IHxQiJAkhMCxXkOg7rtshB069x3Qei8tUukNtnylTuHqFjxFSI0CyAiLWAq0BNA7L2mwUQSuu4lCgttDAGyEKIcQ5c1akQvktRYFTXQJ2EDxnLzZ2DWoPIBsKc3B2Gk2DEaQs0FT9yuTmy4wNjdBiOEZ9Tx8exn6RQKBTuiKnwMd4XkePt+Fhh9igR/X/2zqbHjew6/88599YLyW52t0bSjGacODAGXshINgYMOBtrkY0Bb+W9N1nkS0zrYyQfYXprINvJJpsgq2C0MALDk4FH/5FG6jeS9XLvPee/qCp2NSX5fdxk6/yEEptFNlnFYlfde5/7nEe898F732ZZ1hBRA6BNKYWmaSIzp7quh/yPrT6oJoAYxu2HALhnz575GKMHkNd1PRGRiYjsVVW1F0LYjzFOQwizlNKsDzDf69dNU0qT6XQ6n81m848++uhof39/VhRFqarOOZfleZ4PweY3vbOGYdwyhjoX2g+IDAMjqn32h6zLYGnqBlBYFSwKx11pD8J1h8W2NbjfNjtqnAli7o/dYDPk0RwghmFsNRvnpaGcphKBtLvfOSm766kQ+qBt6ktNMjxncL1Y77wD+tJOytxlWRQlpG26zJAQ4GIAtQEcIzRFSIwgkc79MZTE6t+3H+XvNnXk/liHoev17V7v1uZuDu2GFJFiL7b06epCDO0FDGLuXKO4ytIYQs+7hTrBiKh3fvjO+dE7QFxegIsCPJkARQnJM6S8gOQZKMu6vA/nOvcHEZRdF2TuGIkIkbtA9kSERJ0oldALUUPGx8j1Mez7+NbED8Mwbpo3lfcdt48HMcTaxdtN7wAZAtAbImpUtQXQxhhDSil679P5+bm8ePFCiWirD6gNVhrGLWYIPL937x5XVeWrqspFpMiybFLX9R4RHYjIgYgcpJT2AMwA7BdFsVeW5Z6qTkMIkxhjcXh4uH9wcHBweHh4OJ/Pp5PJpFBV4h7vvXfO2QidYXxrjAtWv3t0To5++EG74PMhCwQxdkuKfSi6rGeKkiqIRyLIFn6Gb3N3bJadG9wg1lnYLjZFj6FTN358mwU4wzCMoSQWgKsB9H4A/ioEvLuGClFXAoupK5elBEYXrO4G4Xe4XmUeGiIQCmgIoBiAEOBigoQWSAmuD1UfxI/hGq7a5ZCsg9HH5a+gnbsTVwP/v1MA6fePh4yRYUCOugVEcOzAwFoAue78IAwePu2Dz8fZH53zxYPzHFyUneOjKMB5jpT5q2wR76GOIcSdmARC4k7sEGLEfnsitBOcgGuix5D1cS3nw4QPwzC2kDdNBBo/9qafjZtHRFRVJaUkTdO0bds2qloR0Tr8PKUUAMTpdBoXi4UA0MePH2+91d0EEMO4xTx58oQePHjAP/zhD9l775bLZea9L9q2nQLYA3DgnDtq2/aOiOyr6n6e5/tlWe4XRTH33k9SSmUIIT88PJwdHR3t7e3tHezv7xdlWeY3vX+G8e6x2b2/RRkfb+Fqpme/DOWvhoGSlECpEz84SR+S3g2aMPpJmutBZ91qGWnoHLwp9NzKYG0vg6ghItfEj82ZbSZ+GIax1YxKRW6KCqrau0AAB0CYEEXhiJH666xz3E1CIAI7B/IOFDNQjNDQ5X5Q7JeUQCF0WV6xD0RPo2D0wbGhV6WvrrV6Rtf0a1fEwX13fceu7SKNBB6g2/YuB6Xbd15PlRg5QYjgBhFoJH6AO+cHegcIsi4AHkUJzbK1+IHB9cEEYYL0OStDlsfa5UFX75eGzx2jnI+N4zM+boZhGNvGptDxtiB0Y3tQVQkhxLquw2q1qler1SqEUBFR5ZyrAbRZloW6riMzJwDp0aNHsu3uD8AEEMO49RwdHdFvf/tbl2WZz7Isq+u6UNUJM8+YeZ5SOmLmO0R0AGA+nU7nd+7cObx3795BURRTZs5SSr4sy3w6nRaz2Sxzzrmb3i/j5njNam8YfzW6AREdHB4iQEqgKKCYQEnAImDtZpAyANcPIoDQRb1u8Sz8NwkbbxNEjO1h0/0hIogx4k1VIbfxe2cYhvG7GDsNtHdCdM6MrkwVq8JxVzKLvQNJlw/CzsHlGTgJKEnv0kzAIICs3Zu9ozP2t9cEkCunB9BNbhgEEIVuTAWhNwogr4Wj82gWMnRd4gq9CCJD7c2+rTDs8+AEUXbdz70AMpT8gnOd2JHnkCLvXR8e4hjqhrJW3Wsl1b6k1eDseN3dIf1WifYuFVjAuWEYu8PQ33qT6DGeMGT9mu0ixiir1ap59erV6vLy8ny5XJ43TXMZY1x672tVbZg5lGW5dn/sgvgBmABiGLeaTz75BE+fPsUXX3xBeZ5zSskRkXfOZSGEIqU0IaIpEe0R0R4z7zvnDiaTycH+/v7R/v7+NM/zjIic934QUZxzzq5S7yDjRso2DyLfVjatw9foe/+3+g+zHwiByigEvZstSsPSD6awKBwUDt2sysENIkNt8y373r6pRNLm39ebauka2wH1YcBZliHPc+R5vj5eIrIWsDaP2+/8mzYMw9gCBvFjOFMNodsJfSZHVzurm3DguBNF2MGDwJ7hFHCiYBU4UWiMYBHIULKyz/8YHJ1IAtIuDJ2GEljosj6Iek+GXrlDGaNz6Xo76VpYerf9V+4W4ivBY+1w6Z88lAJbn65pQz5h7oLQiTrRgxnaiyDqHCjPIN53Yeu+d30AXbA5OrdHFIEoIUkncYjIlcND11s5CmLv9nldpsyuG4ZhbDFv66eMxY/xfevXbBcikqqqas/OzhZnZ2cXl5eX5865hXNumed5JSItgCAi6Tvf+U5qmmYcS7XVmABiGO8Ad+7cwcuXL0lVyTlHRER9bgenlJxzzjPzsGRElBFR7r3Py7IsiqLw3nsmIsv4MABcF0GMvyJDGYhu+mNfyuFdKIQ1Kn0x1AEfZoZKWs8qpT4AfZ0B0g+ecB/mStArEeRmd+camw6P8frx7ZABYmwXzjnkeY7ZbIa6rpFSQggBKaVrnTpmvjYDzo6lYRi7gm7cDgoBoRfsh4wMIjhmKACnXVaIOIB7UYG9h0gCSwaKCdxPZmAA2pe/YtXe9tCV3aLhjWnjvRV9LsfGFV2vnr55rV9neuBKRxDVtfgxfn4n9tAoDL2TTJS6MlhKvBY+wAzpy36J91DvIc4h0VU5q9i7PjoXSF9STId8lU7oWF8z3jYgaNcNwzB2gLe5Pwbnx2ZenrE9iIiGEOJisagvLi5Wi8ViMZ1Ol9PptMqyrBaRlpkjM8vZ2ZksFoudOZAmgBjGLebJkyf42c9+pl9//bVmWZbyPI8AAoCWiOoYYwVglWXZIqXkVdWnlPzFxYVjZl/XtRwdHcnR0dGEiLI3lfMwDOPmuDaYev2RjWXHGaZFrl0gWGeBsGg3i3QIP+8HT1gUHkAa6oeva4h3Aw/bJoK8KStinAkyXm8D59uFcw6z2QwffPABiqLAdDrFq1evcHl5ibZt4Zy7FgI5xo6nYRi7zPiMNrRF1rN70bkvB/9FgoL7DA4mBpyCmUDM3TXauZHTs7t2u5EDY+zyuBaEPrJxUH91XztAhgfXjo5hW7vfW5f36sPHu587sXqzFTUIIV29j94FwgxlhhCBnIMwd4+rQlLsHgPWYkeCQqQrfbV+D9Wr9zYMw7hljIUQc31sP0QkzJy89y0zN334ecXMdVEUdQghTCaT1DSN3L9/Xx8+fLgzB9NGMw3jFvPJJ5/oZ599pmVZiqomVY0iEoiocc7Vqrpi5oWqlkVRcAiBQgi0WCwQQkAIITJznEwm6r0vMDpnqOq6bzHc7wfqiJlp4Cb22/jLsjkL3Ros28XbRZDbw1DmwqnC9Q4PTgmuL33FIutZpCSdGMKqXV1yRV8Ki66JILpV8geuiR2bgYEDMUaEENA0DZqmgXPu2uC6cTN471EUBe7cuQPvPZxzaJoGy+USKaU3Btib8GEYxm1hHJiu6LMsRlkhAlxzZRIIIO2EDwDM3QSHId+D+0kOTISI7nZ4fSgwRHiMkzwAgHEldly5ZXu5ZLiW0rCVQ5mpvg21Fj9oVIpqPJWkSxwR1bXTZXCTvL50+R0iw3sCSfRaxoeMymyZ+GEYxm1iPJFrYBDGmXldMtZ7b23hLYSIlJmTcy445xrvfe2cq5xzVZZljfc+eO9TnudSVdVOXbxMADGMW86LFy/03r17KcaYRCTOZrO2aZo6pbR0zhUxRq+qDCCpaowxtnVd103T1ES0LIpiPpvNKgAT51wGgFSVRYQBkIgwEZGqMjOzc86VZenzPHcWlr7bvGnQztguhlmQQ33r2yiCdOIHIVdFEgGlCIoBHB182yKLAZxiVwqrF0ZYUi+AAAyFA4MhYOrLZWzhQMObBsbHHYeUEuq6xqtXr+C9h4hgb28PZVkiy7Ib2WajYxCiiqKAqiKEAO89VBUxRjDzuvzV24QuwzCMXWZwMxDQ5WT0IogqIJC1KMFEUNLOAdKXtGRiDPGp3J8jmTovB4M6o8XggOxFiqH85/WNGDlFcOUGufr5Kk8DdHW9HVwYxHQlUgyP6VUw+iCA9G/VvTIzkspVQHpfMkskdfclXXu+iPQizNU1YHCgGIZh3AbeNpHLOQfvPZgZ8/kce3t7KIoCNmS0dSiARETBe18zc0VEVZZlVe8GaZ1zqa5r/Z//+R/88pe/vOnt/YMxAcQwbjFEhE8//RRVVelkMkne+xBjZAB1nuccQvD9II2klBpmXjnnlimlhYgsQgiz5XI5e/ny5d5yuSydc7mIOBHxKSUvIk5V/bAuz/NsOp3md+7cmezv75cmgBjGtwdt3FvPj7xlnWgC4FVQAmABiqRAqyAVuMzDNzU4BCB2Igj1zg8eSmFhyA65npeyzUPP40FyIgIzI8aI8/NzqCqWyyUWiwU+/PBDEJEJIFvCWNgQEYgIYoxrgWR4zibmBjEM47agwLpk5YDolYsjaV8ea+3i6ASDcdbV4P4goqsQdCIQDyWw+jbP6LQ5PoNePT5yfozizq8E6F4Joatw9yEfZLO0l47r2ePKxdGVzuLXnSLD54DrzhKMxO+xGGMYhnFbIKK14wPohN+hv7K3t4eDgwMcHR3hzp07mM1msDLr28XgAGHmlogaZq6dcxWAuiiKpneGpP39ffn+97+v//zP/6zHx8c3vdl/EPZNM4zbjT59+lQfPHggR0dHqSgKKoqCptMptW2LvkpVIqJIRJX3fikiizzPpymlWYxxulgsJiIyYeYSQC4ieUopSynlKaUcwPBzNplMyqOjo2mWZSiKgrz31Hcy1uWxRpWxrLlvGH8mwxgDA10f/hb+VQ2DH4UqMiRIEkASoAI0GSi0oBBAKQGpK4Pl+gGKpArXvwavg1S3Wfq4YjMTJISAtm2xWCywXC7RNA3m8zlms9kNbqXxJkQEKaX1slkGwJwfhmHcZlRkPa4vvcAr4/PecD0mWncGBtEioc8I4bWM0U1e6J9LRGu3yCjooxNGaPgdxdr/8VrD6Oq52m/IIHAAb5kc0W+/Ds4WjEQRXOWIjAUO2biGr0WQ9fqr8liGYRi3ibGDbrwuyzLs7+/jwYMHODo6wv7+PoqiMAFk+1iXwCKidnCAFEVRee+bpmmic04A6KNHj3aqU2PfNMO45RwfH+unn34q3/ve9+Ll5aUC0NVqhaIoFIDEGKNzrs3zfFlV1cR7XwKYMPMEQNk0TRlCKFNKpaoWqpqnlAoRKUWkGNaLSLG3tzdh5no+n6eyLCOAVlVZVZ1zjvM89957z11IyI1+Loaxc1z16a+vo+vrbuNfVufi6NSeri3dl5oIAZpiV2IiJegoA4SSdNkfvSNkcIH0v73VLpBxx2FwgKjqOvtDRFAUBaqqQkrppjfXGDFc2wb3x9tEEMCcH4Zh3FLGYsKoxNTVw7SZSb4WObpf7HI2hvJYw5PG4YNDgPkQjD40j2j90/XSVwO68fM4EWS9barXtm8scmC43RA1BjFkLZCs30TXItCuTMAwDMP4cxi3bQdH9LC+LEvM53McHBxgOp2uy8Qa2wMRaT9JOjjnGlVtmLlOKTVZljXOucDMabFY9FFYtDMXNxNADOP2oz//+c/l8ePH+Jd/+RetqkpTSiIiMc/z4L2vASybpsmzLMtVNSeiom3bUkSKXvQoVLUkogJAQUQlgGnvCpn0YsgkpTRtmmZ2cXGxUtW98/PzqYh4IsrLsizm8/lkb2+vzPM8s4D03eBNM5Vt0O4GWVdw0GvlnG41o3DVq1sFVKAqkF74QEqgmMBJABWwaLco1i4QIoB0m6WPjmEAhpmvlcIaBtGHzsSbBtWNm2U4JiklxBgRY1w7QobA+s1sJTufGoZx6xmd58biwLX1w/1h0gJ1IeXah4nT6LHuqXRlhb3mAhkJFd1vjjZk7ETpVBQdl+waiTPrElaj7VtndPUul83nXH9fXHO5GIZh3FZ+3/jAUAaLiOCcQ5Zl5vzYXoYSWIGZGyKqmbnK87wuiqKJMcbVaiWXl5f65MmTm97WPwr7xhnGu4GenJzIyckJVFU+++yz9OLFi3jv3r32yy+/dHfv3nVFUXgi8kTkl8tl7r3P8zzPRSSPMRZZlhVEVIhIGWOchBCm6MSPSUppKiIT59w0xjg7PT1dLJfLGRFNRaRwzpXz+XwGIOV5PlzsHIB1eazhFgCNBoisz7BFjAdbbdD15hhpIHhHJJC30xXh7pwfa/dHAkXpMkCkE0IgI8Go1z+2/Rs8HhwfXCDMvM6TGGZL2eD5djHuAI7D7H/fudOOo2EY7xwjsWF97hyfK4fAc6yfdPWro5cZCxhvPpe+5Yo/OD3Gvzs+R4+cIMO5e50tgtfP59verjAMw/i2GE/W2mQ8gcvGELaf3tEhRBSIqCWimoialFLTtm1omibO5/P0D//wD/Lo0aOdyf8ATAAxjHeJ3olOvYtb05MnT+jhw4d0//59Pjg44PPzc1fXtZtMJn61WmXe+4yZs5RSnmVZkVLKVbWIMZYxxukghvQiyEREJqo6ret6UlXVTFUnIYQyz/MJgP3ZbFZNp9OKiCZElKkq90HqLCLOOee89y7Pc+ecY7NDGsbv4Z0fM+2cINQ7QJBi5wSRXgzpg9AdABpmhvazRxldrfFtdjSNZ0oxM7z3iDGunSF2jtw+huM0hDyq6vr4DbPfgNfdH9v8PTQMw/hrMBaKxyHmbxoue1um1580tPY7BOrNNdfcIhsOFsMwWk10sQAAIABJREFUjHeRzcyP8c/mXt9JlIgSM8deAGkBNFmWtc65MJlMUoxxJw+iCSCG8W6i/UBLP/FJBQB99tln6f79+zyfz+MXX3wRZ7NZe3l5me3v7zdN0zRZlmUxxlxEijzPV6o6lMMqQghljLFMKZW9QDKJMU5SSqWITJbL5f5isTjLsmzeNM0UQBFjLFJKWe8yyYuiKGazWTGfz4uyLMHM7gY/I8PYStatDdq4fdfoi2yrCFQEiBGIERojkDpRhEV7MYQ3Pq9RffAtHrwYOghj94f3fr2YALJ9eO8xnU7x3nvvQURQliXqukZd1+uOn3NXlzbrBBqGYVznD7kuv/XM+dc8p25x+8EwDOOvzVC+97XMp40w9PGtsX1oV5pFmDkACCmlNqXUAgh3794NX3zxRQohCHYs/wMwAcQwDHSuEFXFo0eP5LPPPgMAfPTRR3pxcSH3799Pbdt6Zo4i4kMITZ7nVUopDyFkIpKLSEZEuXMuU9VcREoiKr33BREVRDQJIcxOT0/3m6bZd87NYozTtm1nKaVpjHGaUprO5/O9u3fvSpZl7L1nqwtpGG/mWsDmO4z2weid+0OA2JXC0hh74SOts0AcA0xdICpd6R9bzTgvYiyCDLfjx43tIMsy7O3t4aOPPsJsNsPZ2Rm+/vprvHr1CovFAs65azPkxmH35gIxDMMwDMMwdomxq3nT+THcNwfI7sDMQwms6JxrAbSqGlQ1hBDifD5Pv/nNb3byINroomEYAK6LIOgr6z99+lSKouD5fJ4uLi7is2fPXFEUHGN03ntf17XLssy3bevRZXpkzJx57zMiKlQ1c84VzFyIyHS5XO5VVbWnqjMRmYUQ9lJKeyGE/ZTSXozxwHs/n81mgZknAErvfeacYyIyN4hhjFG8roSogkVAMcKFFj404D4b4/ahXemrpgFVFVAsQWUOtCUQQyeGxNiVwlIFgbogdADUh6fS0Cjf4oHnQfgY538M7g8TQLYP5xyKooD3fn1szs/P1zPiUkrX8ltM9DAMwzAMwzB2mXF7diyCiAhSSkgpXRNBjO0ipSQikmKMqWmaqqqqVQihEpG6D0Jv67qOIYS0Wq3k0aNHsmvuD8AEEMMwRgwiCLohVfr888/13r17cv/+fc7zPBVFwXmeU9M0HGN0k8mETk9PXVmWvFgsHABXlqVLKWXMnInIsBTMXKaUpk3TzFJKMxGZxRj3+2WeUprned5cXFzU0+m0AbAvIvt7e3tTAIX33gQQwxhBo/DQ9TrtxA/f1MibGr6u4GMA6S0UQHrnBzUNsFwA3oPKApjOgNCVw6JeDKLMg6QXDDAErfYvc7N78XsZ54CICLz3axeIDZxvH8Oxcs6hLEsURbEueSUiawfIWPyw42gYhmEYhmHsKmPxY7wMosd4sXbv9iEiqa7rtqqquqqqxWq1WqxWqyrG2BBRKyIBQFwul+n58+fy8OHDbe9CvxETQAzDuMag5KoqHj9+PJzYBAB9/PHH+Oyzz2h/f5/+8z//kz/++GPEGPnLL7+kyWRCBwcHPJlM+PLy0mdZ5pnZM7OPMWYppVJVJ865qYhMRWQaY1zEGC9TSouU0kJVV5eXl8uU0mq1WtUhBOnT0L33Pru5T8UwtpexEYRU4WJAXq1QLBfIVytwaMEp3fBWfguogmIEVyuopK6+VZEDe/tAaIGYoCFCsy4gnZi6wHR2AHVOECaGbPkspGFAfciOGBwE5gDZft5UBmC8jI+fzYYzDMMwDMMwdpE3tWMH18fgAEkprUURY7uIMaaqqupXr16dLxaL08vLy/MQwrJt2zqlFFQ1ElH8+OOP08cff7yT7g/ABBDDMN7CxklNVZUA4NGjR3jy5AkBSIvFggDg2bNnBAA/+9nP6Pnz55xlmRMRV5Ylz2Yzp6q+bdv64uKiJqLKObes63rKzCtmXoQQFsx8qarLpmkWIYQlETVFUchsNiNmFiIS51xGRI4t+dd4x6G3hVioglTgUkQWWri26Upi3dbBVRVQaAEVoCqgdQ1tW2iIQIqd8CFytbADQcEgKFFX+grb6wIZ19IlomtlsMwFsv2MnSDT6RRt265nvr1NvLKSWIZhGIZhGMYuMggc4/5LWZYgIuzv72MymcByXrcPVU0xxma1Wi0vLy8Xi8ViQUSrlFKTZVmrqrGuazk5OdHRJOmdw755hmH8QWwKIm96zvHxMVSVTk5O+PHjx/T06VOeTqd8cXHhQggNgNo5ly2XyyLP86Ku64mqTlV1BmAWQriIMR6GEBbe+7osy1SWpapqSCnF2Wy2l2VZASD/a+yzYewGV3+OBAVEwCmBY4SL8Qa361tG+wB0CAgKbRsgtNDQQkIA9WWwNEQgF8B3YkcXgn49rG8sNGwjQ37E4AIx8WM3ICIURYGDgwOEEOC9R1VVaJoGceNv0/JADMMwDMMwjF1jHGw+Ln2lqsiyDHmeYzab4fDwEEdHR5hMJuvysMZ2oKpJVdve9bFommbRT1xunHOhLMvIzOnx48c76/4ATAAxDOMvTJ8jIgDw8OFD+eyzz3h/fz8dHBzEtm3bpmlcWZZVVVWZ9z7f398v6rqexBin3vvLGOPCe1+partcLuXrr7+OTdO0h4eHqauGxc45ZwKIYQDYSEC/sa3YChRQEWhK0BihMQIxAZIAkS74XAFHhITeRTOIHlsqfgwuAVVdB2cPORLOORss33K895hMJrh37x6KosB0OsWrV69wenq6roM8HNdtFuAMwzAMwzAM43exmf0BAHme4+joCO+//z7u3LmD+XxuAsgWQkRCRNE513jvK+99xcwNM7fOuRhCkBDCTosfAGBlZAzD+ItDRNqfHPXRo0fpl7/8Zfr444/Dj3/84/ZXv/pVU1VVlVJaOucuVfVCRM6yLHtJRN8w84ssy56r6tdN03x1dnb229PT099eXFw8Wy6XL5qmedW27VlVVZdVVa3qum5ijEG6q+xOn5AN40/HvvoKhYpAUuqWGCExQGOCptSVAVu7RtC7QboFWywkDK6AwfExdBhijKiqCqvVCsvlEm3bIt3GrJcdxjmHPM+xt7eHO3furGe9ee9fE69MzDIMwzAMwzB2ifEEnkH8GOd9MDOm0ynu3LmzFkDyPDcBZMvoy80H51ztnKuJqO4FkJBlWSSiVFXVzg84mAPEMIxvjZFCrMfHx8PqBACqyv/93//tfv3rX4e2bdsPPvigPj8/TwASEYmIxE4nSa2qBu99mM/nAqAqiuIghJATUcHMxWw2K/I8z5nZzmnGO8RQW/WGN2NbUIVIQgwBGgIQAihGSIpAb8Meix6E3mGBLjx+G1t0myWRBiFEVRFCwOXlJfI8h6pib2/PZlRtGUQE7z2893DOoWkaFEWxPoZvej5gbhDDMAzDMAxjuxn3U8bih4ggxrh2OQ8lsPb391EUxU1usvF2lJmj9752zlVZllVE1HjvWwAxz3O5d+/ezndQbLDQMIwbgYj08ePH8k//9E/x6OgIy+VSU0orZlYASVVb51yrqktVXa5Wq/Pnz5+fn5+fHwE4bJpm3zk3n0wmB++///7B4eEhee+9zaI13iXe9H1/J/8GtCsNJUk650cI0DaA2nbtAEGKIHVgANyXweItz/5427GMMWK5XOLZs2dYLpc4OjrC/fv3144DY/sY10Yer9sUud60zjAMwzAMwzC2iaFU7+D2GJYY4zUhJMZ4LSfE2D6GElje+zrLspVzbuWcq0UkFEURsyyTs7OznT+AJoAYhnFT6MnJiTx+/BhPnz5N3/3udzXLMmJmFRHx3icRiczcpJSapmlWZ2dnFRGdi8hhVVVHWZa9t7+/H8uyRP+77L13zOyYeV3dxjBuL4MLhPplWLfz7ZM/nj4DRFJCChGIAZQSJAaIJEC1ywFBlwXCTBDVzkIj0pXG2vJB5+E4iwjatl13KlJKyLIMWZYBALIsW7sOjO1i3EF8k9hhwodhGIZhGIaxCwzt2HG7lpnhvUeWZSjLEnmer90gxtagfR6hxBi1aZq2bdtaRCoAFTPXzNwSUQghJBGR7373uzs/wGACiGEYN8rPf/5zOT4+1i+++IK/+93v4sMPP0yr1SqenZ3FPM9jSqkloqaqqlXTNKu2bS9jjJd1XVdlWcYYo+zt7XGWZQyAy46ciBzZSJLxzvCm9sjOt1H+CPpGtwhiCF32RwjgEIDUZ4DIkAHSiR9DCSyIXA9E33KYeT3Tasj9EBFkWbaehbW/v2/lsLaQYebbcPx+13MMwzAMwzAMY9vZnNjjnENZlphMJpjP55jNZsiyzESQLaIvVyZN06SqqkJd13VVVVXTNCsRqZi5BtA454L3PtZ1rZ9//vlNb/afjQkghmHcJAoAx8fHOD4+li+++CLOZjMBIG3bqnNOepEjElEgouCcC8zcxhgFAKqq0hcvXmgIIVZVle7evXvAzPvOOTb9w3i3eNcHThWiChFBShEkXRg6YrqWAcIEsHblr5iwnrW0rYwdAsO2DveZGSKC1WqFZ8+eYbFY4OzsDB999BHu3buHoijMUbBFjDuHg3A1uHoGLAfEMAzDMAzD2FbeVqp1aNcWRYE7d+7g7t27ODw8xNHRESaTiQkgW0Q/kS5dXl4233zzTbVYLC5DCJcppSURrZxzNYA2y7LAzGkymcjR0dHOd05MADEMYxvQ4+NjVVV98uSJPHz4MDVNI0dHRwlALIoiZFnWxBgbZm5ijHWe51FEUgghfPPNN6Gu67ZtW/Heq/eemZmyLMu4w8phGcZtRwHt3R6aEjRGcOrEDyTpnB7oAs+BTgAZTgoE2tryV5sCzTgIHeg6G03TYLFYYLFYoKoq7O3tYT6fW5bEFkFEcM7Be488z5HnOWKMr4la2y7IGYZhGIZhGO8ub+pbjMu65nmOw8NDvP/++7hz5w6m0ynyPDdn+nahMUZZLBbtN998szo/P1/EGC+LolhMJpNlURQVM9eqGpqmSXfu3JFXr17tfAfFBBDDMLYGIlqHFxwfH+s//uM/Stu2iZljVVVBRNrz8/MWQJvnuTRNoyGE1DRNapomqSpPp1Of53lGRG4ymWhRFJmVwzKMd4GhxFVXCktTAmIEYgSNxI/OBdKFoHfKKAGQG93y38f49DV2DQx5IDHGtfhBRFitVogx3uAWG29iKAmwv7+PlBKqqlo7Qd6WBWJiiGEYhmEYhrENDO3SzQk7YwHEe4/ZbIaDgwMcHBwgz/Ob2lzjLQwlsNq2jZeXl83FxcWqbdvV4eHhsiiKlXOucs61RBRUNYUQ9NGjRzvfKTEBxDCMreT4+FgfPnwop6en8fvf/762bZtWq1V0zsWiKNoQQsqyLIpIm2VZIKIYQqCzszNWVarrWg4PDw8ODw/3yrJkm3FgvBu8mwHoikH70HUQepf7ISCVzvWhuhZACACjM32ss0B2ZKB5s2QSM19b3vQc4+ZhZpRliffeew/ee0ynU5yenuLs7AxN05gLxDAMwzAMw9h6xu1V4EoU0XUp4qvJPcb2QkTKzOKci33WR0NEtarWRFQ755qUUjg8PIwvX76Uk5OTm97kPxsTQAzD2FZ0CEg/OjqSe/fuxfPz83BwcBDOz8/D/v5+qus6MXNs2zYRkcQY+fT01NV17dq2BRGhLEvnnCMAYGbqnSA2MmjcQt7xRqZqV+4qBlCMQIrQFLsQdElXLhD0ThAagtABSCeM7NInOIgczAzn3DVXiIkf24dzDnme4+DgAFmWwXu/du40TQMRuVYbedyZBN5cbsAwDMMwDMMw/hpsupWH++N8uyGf0Nqv2w8RqXMuZVkWsixrVbUGUDFzxcx1nuctM4flcpnu378v5gAxDMP4dtHj4+NrJ9pPP/007e3txaZpJMsy9d7HUTksruua67qGiEiWZZrnOaeUZDKZTIqiyL33rs8EMQzjlkAKkAo4Bbi2hjY1pGmAEADpc0B6BwhjrID2zo8dc4AAr4ejO+euuUCM7WKoiTyIHyKCi4uLax1FVb3m4hnu2ww6wzAMwzAM46YZix7D/fEyFj+Gdcb2MXZ/eO9b51zNzDUzr0Sk6p0gLTOHyWSSqqrSJ0+e3PRm/9lYL9kwjJ3i8ePHMplM0nQ6DXme10RUqeqCmc+Z+SUzP1fVZ3Vdf3V6evrVV1999fXz58+/OTs7u2yaplXV7S72bxjGn4CCJSFrW5TVCmW1RFatwCGAUuoa68Abl04E6V9lyxvpm2Ho137ecIDYjKvtZHxshtlyQ4dx8zmbs+wMwzAMwzAM46Z4W/ZHSulam3bcrjW2EyISZo7OudY51zBzTUQ1gEZEWiIKVVWl+XyeLi8v9ZNPPtn5zog5QAzD2CmICJ9++qnu7e1F51y7t7fHIQTvnGNVZREhVdW6riXGKMvlkvqAdJRl6bMs6+pg9cDKYRk7zHjGzTvHMIjcLxABxwivCtQ1tG0hKXaB6CKASl8mSzvHCNC5QvqX24VPcOz42Ky/2995bYDd2F6GDuLQYRwf07EzxMQswzAMwzAM4ybZbI9u9kMHJ/rgSrdMu61D++OhKSURkUREgZkbZq6zLKuccw2ApiiK1nsfvfdptVrJo0ePboWiZQ4QwzB2DR1cIIeHh2G1WrVZlq2yLFsw83me5y+J6HkI4evFYvH1q1evvn758uWL09PTV+fn5+eLxWJZVVUTY0wiYldkY8fZbIjincpBVwAJQAChBSH090W1X7pAdKxD0MeB6K+rn9s+0LzpCBgPjjMRHDPISmBtPeN6yeOZciLyWomzbf9OGoZhGIZhGLeftzk/VBXee0ynU8zncxwcHKAsS3jvrTTvFtH3OaRt27harZrValVXVVWr6so5VwGoATQxxhZAuLy8jOfn5+vyV0S08yMM5gAxDGPnICI9Pj6Wn/3sZ9F7TzFGpJQ0yzINIaQ8z0NKKcUYNcbIq9UKp6enICLUdR0PDw/jwcHBXlmWBdtV2dhB3jSbJomCRSCq6P7dbgbxowGhIUJ0DuI8kGXQPIdkHqnP9nAiQBJoErAqeBBDiF8rh6X6BmVkC3jTMd90DIAIbIPmW8+4NnJK6VqZgDc5Pmz2nGEYhmEYhnFTbGZ/DOuG9XmeY29vDwcHB7h79y7ee+89lGVpfZItQlU1hJAWi0VzcXGxXCwWF8vl8qJpmoWqLp1zFTPXZVk2y+UyTiaTOJlM0ueffy6buby7igkghmHsJMfHxwIADx48wIcffoi9vT1drVZaFEWqqipqB4tIFkLgV69e0Wq1Qh+QTpPJJMvz3APIbnhXDOOPpmtw9j9jMHwoBL37AQQBQYkxtoPQ9Rf5K23tt0cC0BBhSYyWHVKWAUUBKkrAeRAIDgClBEkJLAKIdOIHuHeDSFdNq3ME3+j+/KEMnY+hIzJkgAzihzkHdofNcmbjn9/Z8naGYRiGYRjGVjCeuDNeN7iXvffI8xzvvfcePvjgA7z33nuYTCYoigLOuZvabGMDVUUIIS2Xy+b58+eLy8vLi7quL4loISIrZq4BNCml8OrVq5hlWZpMJvL48WPBrnSSfw8289kwjJ3l+PhYnz17lh48eBBOT0/bLMuqoiiW3vvLsizPi6J45Zx7qaovqqp6fnp6+vVisfimaZqLlJIFohs7zXhwVES7BUBiRusc2ixDlWWonEfNDg11JaJuy5de0e1LQCeCVMSo2GHlPCpmNM4hDNZsEWhK0JSAlIDeEbJ2fozKDW2rcLAZer6+T4BC1y6Qoeausb0QEZxzKMsS8/kc8/kck8kE3nfzkjaFDzuehmEYhmEYxk2w2T8al3AdSmAxM2az2boE1nQ6hffe2rDbhYpIapqmXS6Xq8vLy+VqtVqEEFZEVGVZVhNRm+d5uHfvXrx//768ePFCb9MxNAeIYRi7jB4fH+snn3yCy8tLBaAXFxfqvZeqqmg6nTrnXNa2LfpFRKRk5j0A93B7xoKNdwgdBXcP94fbCHSujzxHKkq4mIAUQTHCS0IhglxGA/87jgJI1IkggdDvf+f64D78nEWQYoRPqSuDJV0pLGIFiQCvVbzS7oW3+AO65gpQdE4XZrC7LoDcpgbrbWIoFXBwcID3338fZVmiqirUdY0Y47ok1uDuGZfIMgzDMAzDMIy/BuPSV5sZdpsiiHMOeZ4jz3PL/thOVFVFVUNKqU4prVR1SUQr51yV53mdUgpVVaWqquSnP/2p/PCHP7w17g/ABBDDMG4BRCSqqicnJwpAJpNJ6tfTZDLh1WqlTdOo916n0+lenudHeZ43zJxueNMN489C+0BvqHTuDwWic4hFCZpOu8faFo4DihigMcCpwm2IKLvKUP5L0JXDSrhqkHNKoJS6jIWUIDHBiYCkD0IXATkGoxMQmPrPk2hrE1Q2XQHXhBDCNQeIiR/bCzOjLEvcuXMHRVFgPp/j1atXePnyJZbL5bojCVzPBNkMvjcMwzAMwzCMb4txf2PcDh2HoDPzNSHE2F6ISJg5MnNLRDURVd77lXOu6t0fsWmadPfu3VslfAyYAGIYxq2AiBSAHB8f64MHD/Tv/u7vaLlcuizLXJ7nJCIkIuSc2xeRo9Vq9YqIClV1zrncOeeIyIpUGjuDAlAaWibU3WeGOIeYeWhRdOWeALAqknZuCFZARZBBwOhrYe5wY1UwFkD6z6HfnySKlGRdBktCBIUEuAQwd2WwiEDUiSDDp0DDa2zZOPNrosdovePu9BVTxHK5xPn5ObIsQ1EUyPPcbOhbBDMjyzIw8/q4tG2Ls7MzANdLYI3Fj/F9wzAMwzAMw/g22cz9GG6Htqz3HpPJ5LVyrsb20YtXQkTBOVczcwVgxcxLZq6897X3Puzv76ehuko/xnZrMF+SYRi3CT0+PpZnz56llFLc399vvPdVWZaLLMsuvPdnIvJquVx+c3Z29vX5+fk3l5eX523b1iJibhBjZ1CgG5xf50AQlKgTQJiRfIboPILzaL1H6xwadqicw4pdl5FBjITdntqhICgIQrQOfl8HwY+s2ZIEEmPvBIldBogoVLrJLUQ0+ji3e6B5swbv1QPrcDucn5/j+fPneP78OS4vL9G2rZVR2jKGjmNZlsjzfB0SmXrX0psCJwdsdp1hGIZhGIbxbbPZHxqCz5kZeZ7j8PAQ9+7dw/3797G/v48sy7a2D/Wu04sZysyRiBoiqgFUAKosyyrnXEtEsa5refTo0a3sbJgAYhjGreP4+Fi//PJLqes6iEgdQqhijEsiulwsFqfPnz9//n//93+//eqrr746PT19Udf1KqUUb3q7DeOPYd0q6ewLnaOBGbp5S4zEjNCLH5fO4ZIdauK1Y2KXUQziTyeEKADpK4OlvpE+lMDSlCBrR0haZ6GMtSTuHSHb5v54E+OsDyaGiqKua7z45gX+78v/wxdffIGXL1+irmsbNN9ixjWUxwLIZrkry3YxDMMwDMMwboL1xDLpHPSTyQT379/H3/zN3+Bv//ZvcXR0hKIorJ26xQwlsIioJaLaOVc551be+5qZm6ZpUghBT05ObnpTvxXMn2QYxm1Ej46OxDmXmqYJItJ471cA3HK5PGfml4vFYppSyrz3RVEUOQCaTqfw3mfM7NiSu4wtZMi8oNF9IupG75kBxyDnoMwg7yDOQR0DznWDqv0scwZQqkD0zSWVdoZ+35UZSg7KBCUGE0FUQYMLZMgBSQmQTgjRPhAd68wMwBEh7YBTYhxGOHQymHk9eL5arhBDhHced+7cuRasbWwfQ2jkdDpF0zRg5mtlsICrY24ZIIZhGIZhGMZfg3F7VETWIggAZFmGvb09HB4e4vDwEM45K4G1xRCR9iWwIjM3zFyllCpVrQDUWZa1McY0nU7lP/7jP/Q29jfs22kYxq3k8ePHAiD++7//O7Iso8ViwW3bctM05zHGIsaYE5HPsixn5iyEoDFGmc1me0VRFMyc3/Q+GMYmBKwH/QFAiUBMADvA9a4P7wDvAecA70A+g8SI5D0E3UCqBxAldQ3YHdY/APTOl27/wa5zgxAhoRN6kghEFUkEHBMQI5AEkE4A6YpoDRkgowFnbPdHM84DIaJ1ACEAhBCgqmiaxsSPLYeI4L3HdDrFnTt3QERYLBZYrVYIIaxn2Q3CxyCOGIZhGIZhGMa3xSB+jBcRQYxx3RYtigKz2QzT6fSGt9b4QxiFoNcAKlVdEdEqy7Iqz/O2KIr48uXLW9txNAHEMIxbCRGpqspPf/rTeHJywlmW1c45yrLsMqWU53mexxiz09PTfLVauaOjo3Tnzh354IMP2DnnvPcmgBhbxTAgP4ggCuoH7QnUOz848xDvQd4BzgPOQ32Eeg8SgWrvIumdD1e1nnZ0QHXsfmG3Lvsl6NwcnfDRBaFL745ASiDpQtFJFaRDBTGCiAJ9Hoiqbv0nM3Z/qCqccxBV+Ezh2ME5D2Z3zSlibBdEtK6hPGSCvHr16lpZrM3jNxa/DMMwDMMwDOMvydhxPBY/hrbpMMFqcIUYO8HgAAnM3DjnqpRS5b1fpZQaVW2Looj379+X4+PjofDErcIEEMMwbi2DCHJ6ehonkwm3bct9jcOciLIYY7ZarfLFYuFFhFXVz2azkpk9ANfDVg7L2AYUAKn24segXRCIGcTcOz48KMtAWQbOcyBGaEqAT4AqiBjaje4DKQEUd0v/6PddmRHZIToH8Rngs27fnYM6B/IeSgzpM04UQEwJNF4GNQjopaRukJlEruer7Eijfhgk984BqmB2EBHUdY3FYok8zzGZTJBlGZxzJohsCYMDZLhNKaFpGpyengLA2r0zdn5YR9MwDMMwDMP4NnhTudVhnXMOzjlMp1NMJhPkeQ4bKtkdiEicc5GZxyHodYyxIaLQNI2EEG5tR8MEkHeb3zv6YZ3s3WDjAmUHbQQR6fHxcQIQ7t27R3meV3meO+cc13XtVqtVVtd1BiBT1WI2m+2paiYibjqd5kVR5CaAGFtDX94Jqp3ooQpwFwBO3ndOj6wXBLIMlOf/tEkyAAAgAElEQVSglMAiawGEiUAKIISr5O8dQpiRvEfwGaLPIM53++o82Puu/Be7q1D43gkiw8yllEAioNS5QKBDCHr3uRARMJSM2qFr4Pg0RcQgAlKKWC4Xa0fB4eEB9vb21h0YYzsYOpN5nqOuaxRFsT4+47IDA5YHYhiGYRiGYXzbjNuhRLR2K8/ncxwcHKAsS+tT7BbKzNE51zBzzcy1qta9IBL29/fTf/3Xfwlu6ZiiCSDvBtdHx1Xx5MmTP7nHfHJyYr3tLeLx48d6fHw8XkWffPLJZmjRrTyB/aEcHx/r8fGxpJTCwcFB3detVACU57lX1TylVCwWi+LLL7+cXF5e0tHREd5///39o6Mj9pbmZWwBQ/krVQUP9/sAcHJdySvyneihRdG5P0Q6B8gwoB9j5xhRBVo3KoG1GygRxHm0xQR1OUGd54jMADGYGdw7QJB5UNbnoDBDgb4cVgKrgkQB6UPS+9PjkAOC3kmhO5abMeRDAID3nfujqmr8v//3NS4uLnF4eIiPPvoIDx4wnPPWWdliVBUppXVpgXEGyBgTPwzDMAzDMIxvi3Fb03uP2WyG+/fv47333sPh4SH29/eR51Y5fBfYCEFvmbkWkTqE0BwcHLR5nsfVaiVPnz69tWOHNqh3e6BhduAgbjx8+JCePn1KAPDgwQMCgKOjIzo5OcGPfvQjAoCvv/76td7z6ekpfec73wEAnJycvPZGp6en9OGHH35Lu9G9/p/7GkdHR7f2j3ZMVVV6cnKCn/zkJ/qb3/wGAPD+++/rycmJfvrppzg9PVUAePbsmX7++ecKAD/4wQ/0ttb0+x0oAPn7v/97vHjxovXeI8aI6XTqmqYpAExTSpPVajVp23YWY8wBZPP5PD84OChveNsNo0NH+RToBvQBdI6OYdC/Fz44RpCk7jmq3cC4c0CMcDGCmQBJEChS1uWDXOevP7D6h7yjMCNlOdJkijiZImU5lLrfdX0WCDkHFAWQ5UCegbPBFdI9Jug/s/HgMfXZKOg+r3W4OHbjRDnsy1AGa7gfY0TbtqiqCiklzOdz3L37noWibzHMDO89yrJEURRIKb02+86ED8MwDMMwDOMvzeaEm6FPlFJCURQoigJHR0drASTLMthc0a1GVVVSSiIiTdu2dYyxVtUaQKOqTQihVdUwm83i//7v/8onn3yyOcH61mDf1N2Hjo+P6fPPP6eTkxPcu3ePfvazn9Gvf/1r2tvbo5/85Cf0q1/9ij/88EPkeU7n5+dUFAUBoMVisZ76m+c5AcDBwQFmsxkBwHw+v/ZGq9WKAODevXsIIWA+n6Oqqr9oL9w5R3fv3v2LvFZKaRfGrf5kQgjqvcd0OtXlcql5nmM6nepisdCiKOSbb77B0dGRTiYTWS6X+otf/EIWi4Wenp7q48eP5Qc/+IH2TpFb/TkNHB8fi6rqv/3bv9HR0REODw/1/PzcEVHpvZ/GGCchhPLi4mJKRGVZlpOU0l5Kaf+mt90wgFHw8WiwW1WhzF3uRea7Af9YrAPPGQRhhvaloagXR1yedWJAniHFAIh07gfg6v8bGGN981terRVmSJZBJjNoUQJZBgbgVQAQHBOSc0CWQbMMmufgvIAbhBBmsPfr3BTtQ9SH6kJjAWHXSkCOXQLDklJCXTd9QLpHXdf9gLoJINsKM6MoCuzv76N3K6JpmrUjhDb+/g3DMAzDMAzjz2WcNTcWQYag864/0eV/zGYz7O3t3dSmGn8gqqoppdS2bds0zappmsVqtVrFGCsRaQC0RNQ65+LFxUV68eLFZiWZW4UJILsJAcAgfHz11Vf8gx/8gJ4+fcrz+Zzu3r3LIQQGwKenp1yWJQOg5XLJRVFQjJGbpmHnHB0dHVHbtuScIwAIIRAAKssSbdsO91EUBfI8v3Z/uVy+9S8jhEBFUWD0mn8QIvIX+2v7NgWQLMt+72s3TfNH/84fQ4wRWZbpcrlUZpayLJWIZDKZiIjoBx98IE3TCAB5//3302KxEAAJgPziF79IX375pZycnEhfHuqdcIQQkX766afyve99L/76179GURQNEa3atr1k5gkzF977qXNukmXZnnPuiIjSTW+3YQBXjdFrAd1DJohzQJaDCwVpH5jMDHgHzTNokwNNAU4JThJ8jMDeHmJoQSJgETCGEkq9FEJdlsT6/dGvfPPWveX+Roj4GxpUY7fF+mkbz6EhzHwo+ZXl8N534o92pawcABkEEO+hWQ7NPFxZgosSblKCy7ILh8881HWOEO3LXg0nwfXJcMcGmLuOyfBxd58gM6/LYjnn1j/f5obtrpPn+XoCSlmWyPMcL1++RFVViDGuj91wLHfpO2oYhmEYhmFsH+t+5uh2WD+UZB0Wa3vuDiKiIYR2sVhcXlxcvFqtVi/ruj5dLpfLPvsjqGq8vLxMP/zhD+Xhw4e3Nv8DMAFkV1gLHkNZqwcPHlDTNPzjH/+YU0osIpznuVNVPjs7c5PJhFNKrmkaR0Tu4uKCATgR4SzLWEQYADdNQ6rKKSUiIkopETPTcrlElmWIMVKWZWv3R0ppuI8YIwGdaLFpe/Peo67r9QjLWNj4XRa5pmlee60/hRgjnHN/ccFh4A8RV8bPd87ppiDyx/w+M7/2ft57DSGoiCgzCzNLXdeS53mKMUoIQQCktm1TlmUxpRSLooj37t1Li8UiHh0dJQDpRz/6kfzrv/6rPHv2TD/55BMBMKi+t/LE9/Of/1xUVS8vL/Xi4qJV1aosy8u2bYuUUsbME+/9hIj2U0rvtW1bN00TmJmdc8TMuxWaYNwqhhwQ9MHeQ+6DOAcuuvqrxAz2DnCuywNpGlDbAiGAU1qHoms/ozwC4P/P3r3suHVldwNfa+29z423IlkXlSzDgGNkIHcPAicBMmjEg5505upH6EFewqXHSD+C9QrfwAECBAhi9MgaJIaRoDuWLakuJA/PZd/WNygeFqtUcstu2yKl9QNKVcVisQ7FIuuc/T9rLeZ1ANJVglyFFVe/7pcBzNUZ6FdbtbkQyzdCje76129r9U1XH+OLIcjV7eC65VdEXM38QNCr63QBSEAE1gpY68tZINpcVsWk6fqNkwTQGGCtIa4GpXcD0nm17evWV3gjwNlC6/+jW9pgbc4FQUTw3kNdN1BVFQBc/j1WSkkgskWMMdDr9SBJLkO+EAIsFguo6xpijOtQ67bHTA5IhRBCCCHE93VbhXEXfoQQwHsPIYR1a1axM6L33i2Xy/Li4uJ8Pp+ftW07Y+al975BRGuMcWmaBgCIb3p3GAlAthwz46NHj6gLPb755hu6f/8+NU1Dbduqtm2VMUalaaryPCfvvY4xamutms/nGhGVUkp3QYhSiqqqUkop8t4rRERmJu89xRgRV698RIRdwOG9X18OcFXREUJYByCb27wKUuDm17qBq865l34N4DIEue3/4rbqkNuCge7yLkDotuWH2vwZr3JbN7fJe78OM75PKPNdAQgzs3MOEDESEccYAyLGGGOs6zporYP3PgBAYGbPzJaIXF3X3hjjlVIuhOCdc/7s7CzkeR7ee++98OjRo3hwcBA//fRTfvDgQQS4rJp41W3eEXz5a8/82WefuTRNm7quK2PMIsaYOOeKEELfe39RluUiTdMlM/fyPDdJkmgiksnB4vW4bcGzq/4AADDm8mpEgIqASAEac3m5tau5IBEgxstB4MwQuh3cVajQDVa//HGXbaJWP/zyetANX6cu9rjalo0A5No2du2lNu7Dy6o+4madyUb40d1ijN1lDIp5tUEMCJeD4Qlh3RLsslJkdf/NZQgCxgAkCUR9OSAdia5+JiJAvLpXu7Jz/7KWSIh0LQCJMUJVVXBxcQFEl+2x+v0+IKIMRN8iSilQSq3nfywWCzDGACLK7BYhhBBCCPGju3lCVRd+3FYB8peur4mfDzNzjNE756rlcjmfzWYz59xCa10rpdosyywAhIuLize68qMjAcj2wpOTE3z48CEBAL333nukLlco9Hw+V845jYg6z3NtrTWrag8dY9Tee6O11jFGrZTSTdMYY4xCRBVCUIioiIgQUTHz5ZrRhhACrc4IXa1XIXbhg1JqHUSswpMuJAGAy8AGYNV+ZfVxZ2MR5trlSqlbQ5FNN2/r2n/USxbou9Dgx3iB7m7r+yw+ICLfdv2b2/sqt3nbbXWL+KsQJMQYIxEFAAje+4CInpl9jNErpSwzW0R0MUanlGqJyBljnFLKJUniEDHs7e358/Pz8Dd/8zcBAMKjR4941SLrjVt1QUT+z//8z2CMcSGEJk3TZQghAYCibduLs7OzQYzxdLFYDIfDYXJ4eNjf29vLtdZKzpYWr0tXlhxXVQoIV22hQOvLgIEuqz9gFQDgatEfVwEIxngZFjBfDgPf7PO6EX7wKni4/Nr1r/M6unjx5bebL4HQDWpfDW7frABhXg8e74IOvrr5dRXGVUSCV5UZvP4HkC/DENrYaY8IAEpdVoB0s1G0uWx7pQ2w0QBaAWh1OVMEESKs+tuubrqbtbIrIUjX/mr12fryywAEIUaGtm3g2bPn0DQNzGYzODo6hDt37sBoNJIAZEt1/Za7g81uP+DmnBchhBBCCCF+iM22Vzffuv3PGCN479f7onJSzm5ARCaioLVujTFLrXUZQqiYuUVEy8xeax3+93//942v/gCQAGQrMTP+9re/pePjY3r33Xfp+fPnuq5rDQAGAEzTNAkiGmZOQggmSZIkhGC896b7XClliqIwxhgDAAYRdYxRAYCiyyRC4WVzd1q1wLoWgsD6ZF289r77eDME2bwc4DLE2OhNvf460VUv+c2v3bz8+4Qgfy78+DFemLuf8aq39V3Xv61i5WW3u3nf+PZVuG6AeVRKhXhZwhMBIGitPQCEGKOLMbq2bdsYY+u9t8aYNsbYKqVaZrZ5nrfM3Fpr3enpqUvT1P33f/+3f/bsmev3+/Ef//Efw+qP4hs3J+Srr76K9+7d88PhsHXO1WVZJoi4aNt2bq29KMvyfLFYjMbjcWaMwSRJlDFGK6UIEbvfc0lDxM9mHX5sDqZjBiSCsPr6ZSByWRnC3gMaDegTwBAAQgDsBkVs9nkFXlV34Drw2Gx31f3sjaX11fvbXxKuAozu2l1w0oUY/GLLK1zdl425IfhdT6+uGmT1s2h1+9TNCVEETApQq/WQ+MvP9SogIQCFwHj5fXEVsuziixyuB7nztf/7rgKEOYB3Di4uzmGxmEPbNkBEsLe3t263JLbPZvjRHYh2iGjdEuvm14QQQgghhPhzNttdbbq5/0lEYIwBrfVLW7GKrcGr6p0YQvDee8vMNQAslVJLrXVFROv5H1VVxSdPnrwVBxISgGwRZsaHDx/iw4cP6cGDBwQA6uzszNR1nWitkxhjaq3NYowZEWXMnGmt0xhjhohJjDGNMSZa63QwGKTT6TTLsixJksTEGBUzqxijQkRCRGLm7g1XlSDIzOtF3e7jVRr8QjP426o9uvBiMwB52YvjywKQl1V7fJ8A5GXVFz/EjSDie13/VUOQ77qtjTM+b7bBAkRkRIzdG1z27Yt4Obg7eO9d27b24uKiquu6CSE0ANAiYh1jbJIkqUMItXOuZuY2hNCEEFoAaM/OztoQgt/b2/OPHj0KqyqQ+CYNTH/8+DEDQBiNRtZa2yRJouu6zpqmKZxzPefcWV3Xw6Zp8jzPldZaMbMqikKnaaoQUapBxM9u83euq9BgAGClLisuuooQipdDvpUGMpeVH13bK1ot9CMzRFwtlL/wg1Y7t3z9CX+9edX1l4LbX7w3vrjRD6ur8OhCkcvL8Cog6cIQxKtv3XgN7j4KzLCu2e02gC7/D7oWYUzqcjZIV/Gxer9qdnp5G6u3XX2BuxxXsp5echkKIYIiAmAG6z3UTQMhBCAiGI32wFonC+dbbrMKpGtFsNn2rLvO5pl78ndJCCGEEEL8OZv7kt0xQbe/6b0HRFzPpRsOhzAcDiHLsu+c6yterxgjhxCic861bVuXZbls27Zk5oVSamGMWSql6hCCJaKQZVm8f//+W3FAKL+1W6Kr+vj1r39NSZKopmlUCMGkaZoqpTIiyr33hVKqj4g9730PEQvvfcHMRQghizGmIYRUKVWMRqPizp07/eFwmGZZZrqwA2B9omzXvgqZGWOMdKOPOG6GF7e1r7otwHhJSPHKX7/5f/Iq/3cvC0F+7EWdVcupH+V2vs/1XxaArKzm9GJXsnYtEKnr2pVl2VhrF23bVt77mpkbrXXFzHUIoSSipXNuaYxZhhCqGOOSiGoiqoio/fbbbx0A+Pfee89ba8Onn34aHz9+/Ea0xfrkk0/44cOH8e///u/9crl0TdPYVThUIWIJAAvv/Xy5XPa//vrrpG1bvVwu6eDgIB+Px1lRFKSUkpUm8bNbL3Li1XBwWC3eUzcYHbo2ObSa+RG7/k5Aq8kaCKt2OnBjxMi1flRXQcvVl26ZR8Ib1R0AcBVxbHy68aWr63ZpSBeE4NUMEF5VgWx87+bNXFZs4HqORxeCMK2qVUitAqGrQIQRIUD3HiByvB6grH7ubtaCbARMiICEQECXIdNqePb1NkqvcVPFn3Vb+4HuciGEEEIIIX5Mm/ueIQQwxkCv14PxeAzT6RQmkwn0+30wq9mTYvvEGKO11l1cXFSLxWJeluVZ27bnbdvOEHFBREsAaPM8t23b+rIs44MHD96KgwsJQF6/9ayPO3fuKABQxhgdQjAxxrSqqoKZi7ZtewDQZ+ZhCGHIzENmHiileojY11oXMcaUmdOiKPq9Xq8/Go2Go9EoK4rCwEbg0f1cgKuQ4bZKje+q3njhTlwlxz9oOeUli2k/OADZ5sWB7xuAvOJ96dphXWtVVVWVJaK6KIpZVVXL1bDvhogqpdQSABbMPAeAedu2pTFm4ZzLELFERL0KQlrvvT06OrLPnz8P/X7fHx8fxwcPHuCjR492elgSIvLJyUnM8xyUUs45ZwGgIaIqhLBUSi2YeV7Xde+bb75JyrLUTdPoJEmo3+9rZpbG+eK16M72BrgKBHgVhjDiZfhB8XIQtoLLWRkbc0MucZc7XF8MXwce65+2fpYzfNfZ5VdzOtbf1337La9jV/M+rj7u5hpcVYBctcFCXN/Y6h6vAqAYoQtRutZavAqHoGvbtaqKYYDLeR+rW+j+v5gZ4mUJxdU8jR0MBzbP4gIEILwagK61AiJaD9nuTl6QaoHt1VXh0iq86h637nkCcBWGxhjlsRRCCCGEED/IzQoQZgatNQwGAzg6OoKDgwPY29uDoigkANliMUZ2zrn5fF49ffp0fnFxcYGIMyKaG2NKrXWVpmljrXVEFPr9fnz48OHr3uyfhQQgrxednJzQ6empStNUv/POOxoATNu2SYwxbdu2iDH2ELEfYxww84CZRyGEESIOjTHDPM8HeZ4PiagAgDSEkEwmk2I4HPaLohjkeZ5mWbZ+depChVc5SP6hYYb4+X1HFYx1zrXD4bAXQqiMMbXWukXEKsa4tNbOrLUDa20PABYhhAIACq11rrVOmbkCgDpN06YsyzbLMtu2rRuPx/6f/umf/D//8z/7jz/+uGu/tZNOTk7iyckJwGUrLBdjtCGERim1VEotYowz731eVZVxzpksy9KmaZIQQrbNQZt4C2xUZABcLurjahEfEQCBAAkuKz5wc67GxvU2vn9dBbhxGWwGAZtVETd/9Te+d+PC9QXrsGYVYqyDkvUcks2ff7WtV9t79Rleuz2EyxySN690FXp0N9W1CYNu3kcXfgBwvHzfVdBca6W1o64FZIiglIIYIyil1n18r4VNYishIqRpCoPBALz3oJQCrfX6ubJZEbL5WEobLCGEEEII8efcnAHSHScQESRJAsPhECaTCezv78NkMoHBYCAzQLYcM0fvfWiapinLspzNZnNjzDzLsoXWuuzaX6Vp6tq2De+++y7/5je/4dWa2BtNApDXB09OTmg4HJrJZGIAIHXOZU3TZMycE1ERQuhba4cAMIgxDgBgEEIYIuKAiIZZlg1Ho9Hw6OholGVZrpRKQgi61+sl/X4/6/f7WZIkhojkcX5LJUmiiqLQh4eH1Ov1irZtrVLKxxjrpmmq09PTftu2/bque8y8IKLRqixukSTJjJmXSqllkiSVUqry3jchhCZJkvbg4KApy7J99OiRZ2YPG1Uou+bk5CT+y7/8S3jy5Ik3xlitdaO1XjLzDAB6IYSEmXUIIYkx5gBQrOas7OT9FW8eXlUydOEGMwPS1Qhx3jhjHADW4cPVBdcDDO7+wY1gYX3hy7xQ+3F17XWJR3cBXQUZdHPU+WXrpq4MYx3zbMwCQcKryhEGAKR1kLKuBum+1FV43NgmvjH0nAHeiDCgu79du6uuguCy8oOAuasAQTl42XJJksBoNIK7d+9CURSwWCygqiqw1oJz1+e3XA8FZRaIEEIIIYS43eZ+Yrff2LW+StMU8jyHwWAAe3t7MJ1OYW9vD/I8l9kfu4EBICBiG2OsY4yl934RQlgQUUlEFQC0AOC11qGu690/AH5F8tv788OTkxO8f/8+LpdLba1NiChrmqZAxIKZ+4jYDyEMmHmktR4x8xAA+iGEPhH1Y4x9IuonSTIYjUajo6Oj0XA4zIwxOsZISimVJIlK01QrpV6YayveHkopKopCE1ExGAxSZg4AwM65tizLumma5OLiIosxZnDZYm1JREsiWgDAkIhKACi99yUiLpRSS0RcImLFzISIMBqN8PPPP+ePPvooroak7GQQ8v/+3/+L9+7dCwcHBz7G2AJAbYxZENEFACQhhNQYkydJMiCiNoQQmDnGGHmjHYmsNonXozv7e2Pxe724vxGMbAYTmy20usuuBRfrMGEjvHiFZ/b6Nq7N93jJdTY+vvrk+vBzANy43tVGcHfTG1Uv3bW6cKS7n+tF4Y1ZIQx81TaL38w081rotaoEuaoAkRZY284YA4PBALTW0Ov14OLiAp4+fQrz+RystQDw4gEsAKyf/0IIIYQQQtx0c9+Rmdfz5rr9z+PjYxiPxzAajSDPc2l7tSMQkRExEpEzxjRa64qIlkqpMoRQMXPtvbdaa5+mafjqq6/i3/7t377uzf5ZSADy88IHDx7Q8fExffPNNwQAiVIqDyH0QgiDGGM/hDBKkmSU5/leURQTY8wEEYchhDyEUHjve9773BiTj8fj3mQy6e/t7Q0Gg0FqjFHd3A4iQiK63u5dvHUQEbXWqigKYma9OhuY27ZNAMAMh0NsmkYTUYKIA6VUrbWulVKV1rpExIVzbt40zcx7fxFjnGutMwBIjDHEzDAYDNAYA19++aWfzWbxq6++iswcdy0E+fDDD/n09DRaa91oNGpjjHWSJAvnXMbMidY6V0oVMcZR0zTVYrFolFJpnueYJInSWr/yzBwhfgqbQ8rjxqLoekYIrIc/rVtCreOEVViy+Tv8smHnf861J/5Lvn1dd4Grbb28A9e3dzOguSWDQYBVVUfX8mv107u5H6v7dfn5VfjR/bzufkP3s96A5+/Ns/43P+7K1btKEKVISti3nFIK0jQFY8x6/oe1dv3ccM6B9x5CCADwYvWHhCBCCCGEEOKm26qIN/chuxasw+Fw3faqmx8oth8RRaWUM8Y0SqkKEZdEtETEChFbY4xFRH9xcbGzrex/CAlAfj744MED+vDDDxVc/r/rVSudXghhFGMchRBGADDWWk+KopgeHR0d9vv9/SRJht77NISQhBDSEEJCRGmv10snk0leFEWWJInRWssrkrhmtSKPSr0wqxuZGcbjMRORGgwGGRHZVUrcrj6uvfeLqqrOT09PT733eYwxXwUCpm1b7PV63LYtjkYj+Pbbb4mI/Pvvv+8fPXoEuxaCnJycwO9+97tYlmXY39+3iFinadqFQyaEkBNR4ZwbnZ+fLwBg0LatWZ0VkRKRUkrJSqJ47V44o6e77OZi6OYC6Y15It3HLyygfo8F1Vd+MtxYqN0MJuCFbViFIl3FxsbA9PXP7MKdG/d5877Gm5e/QSHAzcXvzYCj+1sgwcduuAqsFOR5DswM1logItBaQ1mWUJYleO+vVX3IYyuEEEIIIW5z2+y4GCOEECCEsL7cGLM+EUfsDiKKRBSMMa3WutZaL4mo0lpXSqkaABrvvUvT1B8eHsb/+I//WI/BfNNJAPLzWIcfx8fHuqqqJMuyxHtfWGuHRLTHzBNmHscYp4h40O/3Dw8ODu7u7+8fFkUxijGq1Rsxs0JERUQ6z3OVZZlaVXsI8UqUUpSmqdnf34fBYGCccz0iCqtSuUBEAQBcVVWL8/Pz08Vi0SvLMvPeZ1rrhIhWU4chWmvx6dOnAABNnuc4nU7XLfVXf1x35cWUz8/P4y9+8Quf57ldLpeUpikppTQR6RhjEULoL5fL+ddffz07Pz/vT6fTxHtPSZLoJEnolqBJiK1wLQy5vODmFV78nr/0ZwIAfp8z0F8WRHSDP27c9rXvufF918KbjYAEEIFXg6Nf9r277Gb4tXlZd+bW5qK6nMm1O7TWkOc57O/vQ5qmkKYpMDM0TQNt267nvWySOSBCCCGEEGLTzfBjs/2V9x689xBjXF8udg4rpYLW2qZpWhlj1tUfxphaa90OBgMHAP6jjz4KH3300VsxAB1AApCfw7XwQymVDYfDbubHkIgmbdvuG2OmvV5vvyiKg8lkcrC/v3+4t7d3NBwOp0VR9OHyjP31G1ye3I9KKVRKSesd8b2sWmMRESVpmpobszsYEZmZg9Y6DyGY6XSqENFUVZVaa9MYY+Kco7ZtldbaAIBOkqQEgPp//ud/aDAY2EePHiEAhB2qBOEPP/yQf/nLX4Y//OEP/vDwsDXGQJZlqqoq7b3vW2v7bdvO2rYdNE3TV0pl4/HYxBgzZpbXU7ETfs4n4/f+WT+gZU8XaNwcUXJrC6/N23+D/25ea2W2WgTvhqF3BzhN08DFxQVorcF7D0mSgNYaJKjITToAACAASURBVMjdTkQESZKsHx/vPZydnb0w7+Nl1T9CCCGEEOLttXlM0H3evRHRevj5cDiEfr+/bsEqtl9cCSG4tm2XTdPMnXMLZi611ssYY621bpRSrffe5Xnuv/jii/jRRx/t5PzeH0oW7H5iJycneHx8THC5QJw0TZOHEHrMPPTe73nv90MIB2maHuR5fnh4eHg0mUz2p9PptNfrTdI0HRhj8td9P8SbBVe+6+zf1YBv6vV6MJlMiIjUfD43FxcXpq5rzczovSellGJm1TQNhRCobVsEAMjzHL7++mt+9OgRwGWr/q1/YT05OWFmjv/1X//lkySBfr8PdV1rpVSyGg5fAsCibdtFCKG01vZjjAUABNiB+yfEm+hli7xv+9IvIkKM8dYF8hAClGUJz58/hxgj7O3twd7e3ro6RGyfzRDLGAPGmPXvfvc432xtJjNAhBBCCCHEZsXHzcuZGbTWkGUZ9Pt9mEwmMBqNIMsyOS7YEcwcvfe2qqpquVzOqqq6qKpqHkIokySpmLkJIThE9GmahqdPn8YHDx7syonKPxoJQH5aeP/+fVwul8paa7z3qbW2IKIhM09CCNMQwmEI4VApddjv94+Ojo6ODw8Px8PhcJSmaW6MkcdIvC6otTa9Xq+vtTZJkmgiSpfLpWmaRrdtS0mSkPde68sJ4OC9R601hxBYKRWTJInn5+dwcnLCJycnu/DiyogIn376aXz//fe9tRaePXtmtdY1AFSIuNRal977JREtlVK1UsquWoYJIcRW6A5muo8B4NoZX845mM/n0DQNVFUFzrl1BUiSJK9tu8Wr687iu601wc3WBlIJIoQQQgghNo8HNttcGWNgNBrBnTt3YDqdwnA4hF6vB1rLcuQuCCGEpmnas7Oz+dnZ2el8Pn+OiOcAsCCimojaGKNbLBYBAOJvfvObty78AJAA5KdEJycntFwutbU29d7nIYRe0zQjABgj4hQADtM0PRoMBofj8fhwOp0ejMfj6WAwGPZ6vZ667G0lkat4LVZnmqokSRKllI4xsnMOqqriVfs1UEqh915XVaUAAIhI0WVZidJa471797DX61mAy4EgO/Iiyw8ePIiPHj2C999/3yulXIzRaq0bZq5ijEulVGmMKVeDpFoAeCv/gAghtlO3AL658L3ZAqsbpt00DRhjoN/vg7VW+vzuiJvDKr33oLVeP8abNtscSBAihBBCCPF22az62DxJqmuL282RS9MUhsMhjEajdfgh8wJ3AzPHEIKrqqqazWbz8/Pz8yzL5lrrZZZlNRHZEILP8zwOBoP48OHD173Jr4UEID8NPDk5oeFwaC4uLlIAyJ1z/RDC0Hs/Yeb9GONhURRH/X7/eBV+7E8mk+ne3t6oKIoiSZLsdd8J8dZDIkIAIKUU5HnOzjmcTqdkjNFJkqi6rk3TNEnTNGY1U8QgolFK6RACee+pbVv65S9/2QBAvDFrZGutti+enJzw/fv3nffeAUCDiDURVUqpchWCLJVS7aoCZKvvkxDi7bO56L3Z9zfGCM458N5D0zTQNA2EECQA2SHMvA4/vPfrx7Z7vLuPu4Pcm63QhBBCCCHEm29zfxDg+uyP7mQaAACtNRRFAUVRQJbJcuSOiTFG75yrqqpaLBaLOQDM+/3+whhTMXPLzL4sy/iv//qvu9Kd5Ucncd5PAwGAVm2DMudc31o78t6PQwj7TdMcVFV1SESHvV7v6O7du3feeeedg7t37+4VRZFrqTMTW8gYowaDQXZ4eLh3dHQ03d/fPzTGHHrvD6uqOmqa5o5z7ggADmKM+zHGcZIkgyRJ8uVymXz55Zf6s88+IwBAZt6F01C7PwxBa+2MMTZJkhYRawColVJV1wILpAJECLFlNoOP7vOuQqCb9dGd2aWUurZ4LrZbVwHShR/e+/UBbBdibQZet1UECSGEEEKIN9tmxcfm5zf3I7s3ORlqNyEiE1FYtWdviKhi5goRK0RstNZ2MBh4pVT45JNPdmI+709BFtp/fHhyckJlWZokSVKtdc85NwghjJh5opSa9nq9A6VU1/ZqfzqdjieTybDX6/W01l0LISG2yqodFq5as4H3npfLJXvvkZkVM2OMUVtrFRFRkiTRORcRMQwGA19Vlb937x589tln8PHHH+/Kiy6fn5+z1jru7e25sixbpVSjta4AoIoxVk3T1MvlskFEl2WZNsbQ5X+RrDQJIV6vmy9D3UJ4Vw3QHRA556AsS0jTFIgIkiQBpZSUvW8pRFwPq8zzHNq2vdbPGQBkaKUQQgghxFtus/qja4PbBSCICMYYSJIE8jyHPM9l5sfuYkQMRGSJqAaAioiq1cm7TYzRNU0TyrLkt7X9FYAEID+qk5MT+uKLL/D09FS988472nufOed6McYhAOyFECZJkuwPBoODXq93dHh4eDCdTifD4XBUFEWRZVn6uu+DEC9DK1prveofz3t7e7Cq5lB1XaO1VllrKU1TZmaPiB4AbIzRxhhtVVVweHjIsB4Jsv1VE0+ePOHj4+MQQvDGGBtjbKy1NTNXTdNUs9msMsbUTdM0g8FADYdDk6apUkq9cQHIzTPKhRC7p6sC2Sx9r+saLi4u1u2xhsMhZFkmAciWUkpBmqbQ7/dhNBqtW5o5516o+OkeUxmMLoQQQgjxdtnc97s5+0MpBUmSQFEUMvdjx21WgCilGkSsAKAmojrLsqaua1dVVTw/P3+rF3IkAPlx4MnJCX799dfqV7/6FSmlzMXFRWaMKZxzwxDCnvd+3zl3OJlM7hweHh6/8847x/v7+5PRaLQ3GAwyrbWcqid2htZaDQaDjIio1+upfr+ffPPNN2o2m+mmaZRSionIhxC81rr13rer91DXNX/++ef80UcfMexAFcj9+/e77QxE5IioJaLGOVedn5+XZVnOv/nmm4vJZJIeHx8jEfWUUvQmn30rQYgQu+e2ahAiAuccnJ+fQ1mWcHFxAQcHB3Dv3r31WWFi+xhjoNfrwd27dyHPcxiNRvDs2TO4uLiApmnWB66bra8k9BBCCCGEeDttVn50Mz+MMTCZTODw8BAmk8k6BHmT1zHeYIyIXQBSE9GSmasYY+29b0MIjojCkydP3tr5HwASgPwouvCj1+vpuq61UipNkqTw3vdDCKMkScZZlk0R8WB/f/9gf39///DwcDKZTIbdzA+llMSsYmesWlyZ1UI/IiJVVcUhhK60wwFA45xrlVIVADRVVbVFUUAIga21XRXI1g9EBwBYLpfc6/UCEbkYoyWiJoRQV1VVO+cqIlq2bVvleZ4dHR1lMcatv09CiLfHbYvgXRWI9x7atl3PkNBaw/7+PvT7/de81eJliGjdrqyb6VKWJczncwghXDtwvW3wpRBCCCGEeHNt7vNv7vt1+/tdlXCe5zCdTmE6nUKe55AkiVSA7I4YY+QYY7DWttbaxntfI2K1aoNVW2vbEIIdDAauruvwxRdf7MRJyD8VCUD+QicnJwQAdPfuXTWZTIy1NkHEnJl73vsBIo601tNer7ff7/cPj46ODvb396eTyWTY7/d7aZpmr/s+CPF9de2wjDEaAIiZcTQarQMN55x1zlXe+5qZl9baJk3T1nvPRBQnk0n88ssv4wcffLD1s0AeP37M9+/fj+PxOFRV5cuytADQxhibpmnqxWJRxRirJEmaw8ND570PLCtMQogt0h0AvWwmiLUW6roGRIThcAjWWlko32Jd8GGMWT9+SZKs2111PZ5vm/kij6sQQgghxJvrtn29rvqjO/mpOyZIkgT6/T70+33IMlma3CUhBA4h+KZpbNM0dVVVlbW2ijFWzFyvhp83zjk7GAz8H//4x/jo0aO3+kBAApC/DH7xxRf4q1/9StV1bQAg1VrnRNRvmmYUYxwDwLQoiv07d+4c3blz5+50Oj0cjUZ7WZZlSmrLxBtAKUVFUZiDg4NenuexKIp4cXFRz+fzsq7r2ntfJ0liich67znLshBCCG3bxs8//zzuQhXI+++/z//3f/8XQwgeEV2M0QJACwANEbWIaLXWTinliShu+/35PqRlihBvjtvaIHUL5ES0Hnwuz/vdsdnS4GbIcVvfZyGEEEII8ebqToC5+da1v+paYHnvwXsv+4g7KsYYmqaxs9lsvlgszsuyPK3r+sI5V3YzQACg9d67s7Oz8OTJk7e6+gMAQGqb/gLMDOPxmNq21SGEJMaYxxgHVVXtWWsnzrl97/2+1nq/3+8fHB0dHRwcHEz29vYGaZomRCQBiNh5WmtMksSMRqN8MpkMDg8PR+PxeNzv9/fTND0wxhxorfe99xPn3HCxWPTats1ijGY6nSpYVZC87vvxMp988gkvFgt+5513AgCEJEksIrYhhEYptX4zxrTGGE9E8XVvsxBC3HQz/OhK37vAQykFiAjee2iaBqqqgqqqwDkHMcrL2rbqHrskScAYA8YYUEq9EHrcVgUkB7xCCCGEEG+Wm/v8m/uEiAhaazDGrPcd5cSn3cHMHEII1lpf17Wtqmp5fn5+fnZ29vzs7Oz5fD6/cM4tsixbElHTNI2NMfpnz55FANj67is/NakA+Qs8fPgQf/GLX1BVVZqZkxBC1rZtn5lH3vtxCGGMiGMAGBtjRkVRjHq9Xl/aXok3CSKS1houR9koJqLYtm3rnGuJyCNii4jWOdcAgNVat8vl0hKRPz4+dgAQ4PK1HLa5cuKrr75iY0zw3vsQglVKdRUgDRE1xhirtXaIuPUVLUKIt8/Nxe7Nz7sKkBgjOOdgPp+vewD3+31IkgSSJPm5N1m8AiICrTXkeQ6DwQBCCNeqQWKMLwRfALfPhRFCCCGEELuta4kKAC9UBSul1uHHcDiEPM8lBNkhMcbonAtt27rlclmXZVnO5/OLxWJxvlwuzxBxBgClMaZm5mYwGFhrrQeA8DYPP+9IAPIXuH//Pv7pT3+iGKMmonS5XPaYeRhCmHjvp23bTohor2magXMujzGqbT7TXYi/FBGpNE3Tvb29kTEm1nWNy+XSV1Xlm6ZpiKhZ9SNse72ee/r0qfvqq6/iP/zDPzBcBiFbZ7VAFB8/fhy+/PLLgIhOKWW11u2q8qNeBSDNqg1WkABECLELusXvroogxgjz+RxijFCWJZRlCe+88w6MRiMJQLZUF34cHh6CMQb6/T7MZjNYLBZgrYUY47Vh6Z3NihCpBBFCCCGE2H03q3+72XDdyTFZlsFoNILxeAzj8RgmkwnkeQ7SnX83eO/jcrlsz87O6rIsZ4vF4rxpmlNmPtVanyPiHBGXSZLURGSZ2ed5Hn7zm9+89dUfABKA/GDMjL///e9pPp8rY0xirc2YuRdCGDHzmJknxpiJ1nrPGDNAxBwu/78lABFvrNVgdNPv9/vGGMiyDBHRhRCctbaOMVYAsETEuq7rNk3TdjKZeLgMP7b1RZkBAP7t3/6NASAopTwzO2ZuiaglokZrXSulGlj1WPTeB6VUICLsvN67IIR4222e7b9ZBt/N/uj6Anetr5qmAe89jEYj6PV6r3nrxcsopSDLMhiPx+tKHWYG59y6r/NmJYgEH0IIIYQQb6bN/buuCqTbxyciSJIExuMx3LlzByaTCfR6PUjTFIhkOsIuCCHEuq7d+fn58uLiYl6W5bnW+hQRz9I0PSei+WrNrVVK2RCC//jjj9+oGbV/CQlAfoBVFQcmSaIAQDNzAgBZCKHvvd8DgGmapvtJkuwPBoPJ/v7+cDAYFFprg4jyyiLeWESERKSVUlophVprjDE6Zg4A0Hjvl8w8994vEbFp27bRWvvPP/88LBaLrR6IPh6P4zfffBMAwCOiIyJrjGlCCLUxpooxLpumWc7n8yUi5r1ej/I816vWYDsZgNwcnCaE2G23zYHYnAUSQgBrLTRNAzFGMMZA27brYYli+3QHs107A6UUOOfWj1ld19faYnUHuPKaLoQQQgjxZuqO37t9wO5EGKUUFEWxrv5IkkTaX+0QZo7OOVuWZdUNPx8Oh8+LonheFMUpM8+01iUA1Mvl0v3VX/2VR0QZ5rgiAcgP9Nlnn5FSSiVJYqy1qXOucM71QwgjY8w4y7Lp4eHh5M6dO5ODg4Ph/v5+URSF3tWFUCFeEQKsh7KqJEmyXq83JqKY53lT1/VsuVye1XU9d85VSqkqxmj7/b7L85xge9tgMTPH3//+93E+n4c0TZ1SysYYW2NMrZRatm1bnp6ezr33s/39/WQymcD+/n7R6/VQKfVGBJ8ShAix+26b+dBVgYQQroUkckC0O7qD2jzPYTKZABFBnudwdnYGs9kMrLXXKn82+0NLNYgQQgghxJthc+5HVwXsvX9h32/zvdgNiBiVUl4p1Wqtl0qpORFdpGl6lqbpBQAsiKhGRGuM8X/4wx9kB3+DBCDfHwIAHh4e0rNnz3SWZYm1NkPEQik1IKJRmqbjwWAwOTw8HL/33nujyWTS7/V6aZZlO3smuBDfFyIqIkqzLEOtNaRpWiPis7quR977c0Qsm6bJkiRprbU2z3MLl8+vrXyRRkT49NNPY5Ik4fz8PBCRA4A2SZIaESvnXHl6ejq/uLi4aJomZWbd7/dNlmXSUFMIsTVedqDTLaDffBO7o6sGGY1GkKYpGGPAOQdVVUHbtusDYWmDJYQQQgjx5tncr9uc/dHNguvey4lOO4uVUj5JkiZJkipN07nW+iJJkoter3cRYyy9900Iwc1ms3BwcCDVHxskAPmemBl+//vfqzzPzXK5TAEgJ6Ke1rqfpukwTdO9fr8/2d/fHx8cHIym02lvNBplSZJoGQUg3iaIiEopRUQZEUVmHmqth4g4iDH2Y4y9JEmW1tpmNBq1y+VSf/bZZ90skG3Ejx8/5slkwtba0Ov1vNbaMnPDzKW1dtG27cI5t0iSpDcajXLnXC/GKKtLQoitcrMSAACuDcpWSsnB0Q4iIjDGrMMra+26tUF3BuDmPJBNEoYIIYQQQrwZNjs3KKUgTVNI0xSGwyHkeQ5aa9nH30FEFBHRa60brfVSa12maTojornWekFElda6YWZXVVV49uyZ7NxveCPasvycfvvb31KSJMpamwJAwcwDZh4aY/am0+nk/fffn/71X//1/gcffDC+c+fOoN/vp0mSrNaBCUGGoIu3BwIArSpBNCKmIYQihNCPMQ5ijAPnXB8Airqu06Io1GAw2OrnyMnJCadpGgeDQej1eg4R2yzLKmPMYjVwam6tXXjvqxhjCwAetjfQEUK8pTYrALrQA+ByAV1rDVrr9SL65tfF9usCrO4xREQIIazfutYHALe3QxNCCCGEENvvZSeubLa+IiJI0xSm0yncu3cP3nnnHZhMJjL4fEetWmA5pVRtjCm11jOl1ExrPd/b21uMx+NKKWVns5kfDAbh8ePHEoBskN/472k8HlNVVTqEkNZ13Qsh9EMIQ2PMaDQaje7evTt+77339u7evTuaTqd5mqZ6FXwI8dZiZowxqhhjEkIonHMDZu4TUWGtza21aV3XKs/zrX+uPHnyhLXWMcYY0jR1zNwkSbIkolIpVRLRkohqpZQlorCtQ92FEG+3zTP+uxkgXSCy+Xl3AHVz8Vzshs2QY7MKBODF/s9S8SOEEEIIsRs299luzurs9vkAANI0hclkAsfHx3D37l3Y29uTAGS3MADEGGNkZo+Irda6IqIlIpbMXCqlysFgUFVV1c7nc/f06dPw0UcfxU8++UTWojbIb/z3g3fv3lXz+dxUVZU3TdN3zg1jjMMY44iIRnmeD0ajUW84HOZ5nidaa5K+V0IAMrMKIaTOuSLGWDjnes65wjmXLZfLxFqrnj59SicnJ9v8fOH79+9zkiQxhBAQ0fX7/UZrXSmllkS0BICKiBpEtAAQJQARQmybmwvg3SJ596aUAmYG7z0sFguYzWYwm82gaRpwzr3OTRevCBFBaw15nsNgMIB+vw9Zlq3numwGId31AaQqRAghhBBiF9ysANms/Ogqf7v5H3mew3A4hNFoJC2wdkwIITrnXNM0dVVVy6ZpSu99CQDdybeVtbax1rZpmtqiKHye5wEAWNairpMZIK8GAQBPTk4IAHTbtmmMsQCAvvd+GEIYhRCG3vsBMxdE1LW9kumhQqwwc1cBknnvC2YuYoy59z4zxhjvvUrTtPsrvLXD0B8/fsz379+PVVUFY4xjZqu1rpVSFSJWRFQRUauUckQUYEvvhxDi7XZzGDbA1RwQIgJmhrqu4fnz5xBCgLZtYTKZwHA4BGPM69x08QoQEYwxMBqNwDkHxhgoyxKqqgJr7fo63fuboZgQQgghhNhONyt8u/24LgDZrN4OIYBSCowxkCSJVH7smBijr+u6KctyWVXVxXK5PK+qah5CKJVSFTM3xpi2qio3n8/D06dP48cffxxB1qFeIAHIn4cPHjyg8XhMAKDSNDUhhJSZC+/9wDk38t6PnHMja23fe5/GGBUzyxGkECvMjMxMIQTjvc9jjDki5t77XCmVIqJZLpfae0/3799HZuZtXYQ5OTnhf/mXf2GtdUzT1DOzJaJGa10xc83MDSK2iOhXQ6rkD48QYqvcXPjefL3t2mCFEGC5XIK1FhaLBZRlCUQEWZZBURSva9PFK1JKQZZlMJ1OIU1T6Pf78Pz5c/j222/BOQchhBdaXt2sApGh6EIIIYQQ2+Vl+2mbwYf3fv2+u1zsJu+9r6qqevbs2dl8Pn++XC5PQwgzuKwAqRGxnc/n7u/+7u/co0eP+PHjx/zxxx9L9cctJAD5buvwo9fr6TzPtfc+Y+airuuBUmovTdPJcDjcHwwG+9PpdJzneaG11rDFg5yF+LmtZoCQ9z6JMWYxxoKZC2bOmTn13hutNRERPn78eOufO+PxOH7zzTeh1+uFoigsM9ez2axeBSD1qgLEwuUAdPnDI4TYOrctbm/OAOkOmtq2BWYGYww0TQMhhNewteL76ipAiAiMMaC1BmYG5xwopaCu6/UZgzd7RnfvpR2WEEIIIcT2uFnBvTnfrav4iDGCUgqKooCiKGA0Gl1rgyp2SwjBO+fqsixns9nsbLlcniZJcqG1XiRJskTEttfrOQCIDx48YETkk5OT173ZW0kCkO+GH374IQKAqqpK93q95Pz8PLPWFt77gdZ6lGXZ5OjoaDqdTqcHBwd7/X6/p5QyMvdDiCuICKvKKL2aA9JVgGRa6xQRE0RUdV3T8fExPnz4sHv+bGN4wI8fP+bj4+M4Go08IjpmbhGxjTE2IYSGiCwiekSUUy2EEFvpZvXH5gwQIlqfKdYFIV3VgFQF7I7NgfbdTJcuAOnaYXWPa+dmOywJQYQQQgghts9mVUcXfHjv13PgBoMB7O3tXWthK/t0OynGGK33fmmtnTdNM1dKLZRSy1X7KzubzYKsPf15EoC8HD548ABPT0/VdDrVRVEYZk6VUnmMsRdCGCilxoPBYHrv3r2Do6Ojg8lkMi2KIsuyzBCRvLIIsXLZ0QoxhGBCCEmMMUXEjJmzEEJKRAYR1eHhIR4eHsJXX321tTNAOk+ePOF333035Hnu6rq2McbGe98wc8vM6wBESg+FENvqZSFIt2jenUGmtQal1Astk8RuQERIkmR98FsUBZyenq7bJDjnXtrySh5vIYQQQojtcNvJKZvDz733kCQJZFkGBwcHcOfOHZhOp9Dr9SDLMtmv20FEFJRSzhhTGWOWxpiFUqpUSlV5ntcA4JMkkRL9VyDTb77Dhx9+iFprAgBdFEVS13UeYyxijP3VwPMBEQ3yPB+ORqPB3t5eURRFopRSUgEixJXVoplK0zTp9XpFv9/v5XmeK6UyZk4AQDOzquua8jxHgNvbs2yLk5MTBoD4xz/+MT579iycn5/7tm1djNExs7XW2uVyaefzeTubzexyuXTOuRBC2N47JYR4K93cXemqBhDxWvjRXS52TxdqZVkGg8EA+v0+FEWxboXQtUzYbIe1WREkhBBCCCG2w+ZJK93+W7ffnuc5DAYDmEwmMJ1OYTqdwng8hqIowBjzmrdcvCKOMUbnnG+apm2apnHOLZm5JKIFEZVa69IYUymlWkT0dV3LOtMrkAqQlzg5OUEAoNFopJIkMdbatCiKoizLgXNuaK0dhBD6zNxPkqTIsixP0zQlWR0Q4gWIiMYY3ev1svF43DPGNNbavnMuizEm1loDAHowGNDTp0/p4OAgwuUcnW19IedPPvkEHj16FAEgNE3j27b1MUYXY3TL5dKenp42Sql6PB7Xk8kkH41GSZ7noKT5phBiC91c/O52Z7oqkC4EkQXx3dQ9hsYYqKrq2kwQ7/210EsIIYQQQmy3zRCkq/YtigL29vZgPB7DwcEBjEYj6PV6r3lLxfexmucS6rp2TdO0VVUt5vP5wns/jzEutNYLRCyJqELEBhH94eGhtL96BRKAfIfJZIJnZ2dkrTVJkqTOuR4A9GOMA+9931pbOOdS771mZlkREOIliAiTJFGj0ShL05SXy6Uty7I3m82yqqqSEIJOkoTatqUPPvgA7927t/XPJ0SEk5MTPj4+ZgAI3vvQtm2IMYbz83NrrW3Oz88X+/v7/ePj45yIUGuNSZLI6pIQYiut5jWtzyTrFsS7N6kIeDN080CstWCthbZtQWsNWut1+NUFYJtD0eWxF0IIIYR4PTY7ZHQfd/P5tNZQFAXcvXsXJpMJ7O3twWAwgCRJXtfmih+OnXOhqqrm7OxsMZ/PZ1VVXTRNMw8hzJVSpTGm0lrXWZbZGGNYLBbbeuLwVpEA5CW++OILvHfvHh0eHqqmabT3Pg0hFN77Xgih773vWWvztm1T55yOMUrlhxAvh0oplec5aq151foqrevatG2rAUAxs0qShM7Ozmg+n+P9+/dxNTtkW1/MGQDwyZMnPBwOGREjEYUYY1gul95a285ms8Z73+R53h4dHaXSAksIse02B6B3i+GrM5GgrmuYz+eglIIkSdaL5mK3EBEYYyBNU0jTFJxzAADr/tHdY969QpdUZgAAIABJREFUB5BZIEIIIYQQr8N3zfzo5rkZY9bz3sbjMYzHY9lP31FdBYhzrlkul4uyLC+qqrqIMc4BoFRKLUMINRG1iOhGo1H46quvZJ3pFcii/Us8e/YMR6MRtm2rEFE755IYY+6973nvezHGPISQOueSEIKSChAhXg4RUSlFxhidZZnJ89zkeW6IyACAVpfIe6+Oj48xSRL87LPPtv45dXJywl988QVrreNyuYzMHGOMoW1bP5/P3fPnz+35+XlblqVzzgXe5sEmQgix0rVD6t6YGdq2hdlsBqenp/D8+XMoy3K9cC52i1IK0jSFwWAAw+EQ+v3+ui90VwEEANcqgSQAEUIIIYT4ed2s+th868KPrgqEiCBNU+j1etDr9SBNU2ltupsYEX0IobXWLpqmmTVNMwshzBGx1FpXSqlaa90SkZvNZvHx48eyzvQKJA58iY8//hiePn1KxhiVpqlBxJSZ81UFSM85V1hrsxCCCSHoGCNJCCLEK0NmJmZWMUYdQtBaa6W1ptlsRlmW0WAwiKvrwTZXgXz44Yd8dnbGzBxDCAERAxH5GGMgIk9E3WVxi++HEEJcO8jarP7w3kNZltA0DZydncF4PIZ33313PVhbFsd3S5qmMJlMQGsNo9EInj17Bs+ePYOqqsBauz6w3qwAAbg+dFMIIYQQQvx0bu5zdfvbm5UfMUZwzq2DEPFmQMSQJEmdZdk8TdMLZj4nohkALJIkqYiottbaoij8Bx98ED/66CM+OTl53Zu99SQA+Q79fh+ZGUMIioiMcy7z3mcxxiyEkFhrTVVVejab0fn5OWRZxlmWQZIkXa9sWREQ4gZm7p5XFGNUMUYVQlAxRnLOERHht99+i3me78Tz5+TkhH/3u9/xYDDgGCMTUWTmiIghXvaRiYgo4YcQYuvdLK/vzvwPIaxDkKqqIIQA4/EYJpOJzIbYQcYYQEQwxqyHoVtrAeAq+OpsVoNsXiaPuRBCCCHET+Nl+1qbg8+763QtTdM0Ba31tf04sTM4xnjZTiQE65yrY4ylUmpmjLmIMc4QsQSAipkbY4wdjUbuT3/6U/jggw9krekVSQDyEl9//TWmaYrMTMYYxcyamdMYYxpCSGOMibVWl2Wpvv32WyyKAgEAJpMJD4dDzPNcDg6FeInVohoCAK0qQYiZFREhEeHdu3fh/PwcHj16hA8ePNj2F3P+9a9/Hf/93/89MnP03kcAiCGEiIgBACIAcHdGrRBCbLPbzvLvzi5bLpdgrQWlFDRNI2ea7ahuqH2apgAA8P/Zu5ffyK7jcPx13vf2u9nkPKRJbClCENCBN/ImuxHgVfbjddbJHyHqz4hXwXep2RrI0tbWgAMESQhkIxuxftLMkOzHfZ97HvVbsO9VD83RcySyOfUx2qQ4HE6T3X15TtWpKu89NE3TD713zr20sd7dhFPygxBCCCHkx9etyXbXaFprMMbAdDrth55TAmQvYYwxOOdcXdd10zSFtTYDgLUxZh1jzDjnBQBUnPMmhOAGg4H/+c9/Hij58c1RAuRrKKUYY6xv1RNjVCEEHWNUVVWJGCP/3//9X7bZbHC1WsV3332X/+QnP6ELDyFfYdsurmuDxbcY55xVVcXTNGXHx8dwfHx803f1G3n69Cn8zd/8DTrnMMaI3nvknMedChD6pUQI2RvdpirG2FeBCCH6YYpSyq7S9abvKvmetNYwHo8BAGAwGMB6vYbVagVVVYG19qXPpSQ+IYQQQsgPb/cAynXr7W7w+Wg0gqOjo74yezKZ9HPdyP4IIYBzzud5Xq3X63VZlufOubMY4zkArJIkyQCgZIw11loHAH6z2VCc6VuiBMhXsNayEAIXQnAhhEBEGWNU25kFom1bUdc1q+uaZVkG1loYDAZweHgIs9nspu8+Ibda1woLLmekM8YY897zyWQCFxcXLM9z9t5779303fzGNpsNaK1xK24HnkfGGG7f725767qT4XQamJC7ZffUf4dzDpxzEEL07zvnoGkaqKqqb6VEgxb3j5QShsMhaK1BKQVCCKiqqq/wedVjSvNACCGEEEJev6uJj912pDFG8N6Dcw601n388ejoCGazWb+eI3sHvfe+qqrq/Px8XRTFeYzxPE3TC2PMSim1CSGUiNhVf4RPP/003vSd3jeUAHmF1WrFhsMhAwAmpeQhBA4AYjuzQCKicM7xtm15URRQ1zUYYyDLMmjbFi4PfhNCvkqMsW+DxTnnSZJAURQMAOCzzz5jn332GXv8+PEN38uv97Of/QzX6zVyzjHG2CU8IiL2FSD7mJ3vFl3XnTyhll6E3F1XE5u7VSBCCEBEqOsasizrT591rT+p+nW/cM77vtHdLJBu49xttDnn/XOgW9/S9Z8QQggh5PX7qn13N/g8hACICFJKGI1GMJlMYDKZ3MTdJa8Hxhi9974piiLPsmwDAGsp5TpN040xJhdCVHVdW0T06/WaAs7fASVAvqEYI2OXR7kZIrIYY3d76YJEG0JC3lzWWrgsFvvyQrB9d+8vDJTwIOTN1SU2lFKAiGCthfPzc3DOQVVVcO/ePVgsFiAlLSv3HSKC976/SSn75AciAuecDvkQQgghhPwIuj14l/jw3kPbtuCcA+99nwghew8ZY5Ex5qSUNee8RMScMZYxxnLGWBVjtADg7t27551z8fe//z098N8SHdP7GiEEFmPsEx9dy57trWvjQ8FBQt5w6/UahBD9RWCnEmSvLwxXr22771PrK0Lupt32RrvVH10lgPceNpsNPH/+HJ49ewabzQbatqWh6HfAbqXPdXNeqO0hIYQQQsgPY3cNvhtn3F2L77ae7dbmZC8hIsYYY/DehxCCQ0TLOa+EECUAFIiYI2IphOgTIMvlMuR5jh9++OFex5luAh3V+4a2iQ6+vfVJke2fUQKEkDec1rq/AHQtr2KMCJfZ/L1sgUUIId2mq9twdX2HuzkRUkqo6xq89zd9V8n31D3Gg8EAhsMhhBDAe9+3WrjaFvFqcpw24IQQQggh393uLL7uxjkHKWVfib0dmN23vtJa0xy+PbTNfoS2bb21tq6qqmyapogx5gCQCyHyGGMeQiidc/VoNLKr1crdu3cvHh8fUzn2d0AJkG9gO6fgq9COj5A33GAwYNte6UinoAkhd0W3CeuC3t0w9N2B6BT4vhuEEDAYDODevXtgjIE0TWGz2UBZluCcu3Y2DCU+CCGEEEK+v93q693/VkrBeDyG6XQKxhgAAIgxgtYaJpMJjMdjGny+hxAR27b1WZaVWZblRVGs6rpeWWszAMgZYyVjrAKAejQa2TRNXYwxvPfeewG2h2xv+FvYO5QA+QauC2huN3204yPke+Cc4+VoHXxpbsZdIYRAzvnet8EihLx5rgtq754u64Zjc87702je+z5BQkHx/SOlhDRN4ejoCIwxoLUGAOjngQD8ZaXH1SRIjJEee0IIIYSQ7+Bq9QfA5fpsOBzC0dERTCaTvhKEcw5aa0jTlObw7aEYI7Zt64qiqJbL5Waz2Szbtl3HGDPGWME5L7ftsBqtdbtarcKLFy/ie++9R7Gl74heJd/QNkj70se2gU0ACm4S8p3RMFVCCLmddk+i7bbCijH2FSAxRmiaBrIsAykljMdj0FqDlBI4p1Fz+6R7zHYHn1troW3bfvBmN4SzS3J0z4GrpxYJIYQQQsjX2z1I0iU+Yoz9eosx1ld7zOdz0Fr3H+/W5rT+2kuIiL5t27osyyzLsk2McaOUyqSUhZSyYoxZ51z76NEj9/TpUzw9PcXHjx9T9cd3RAmQr7E71Hj7JEPOeXeq+6ULD110CPluugqQpmlgNBoBAMCjR49wn7Pb21PR3awgujgQQvbO1TkPHSFEn7x2zsFyuYQYI9R1DYeHh3BwcACDwYASIHuoq+pJkgQQEbz3IISANE1hvV5DURR9pU9X/bO7/r2DxZyEEEIIIa/ddYmP3fe7tfbuISQpZd8Gi+w9ZIx5AKgRMQeANSKupZSZlLLgnNdKqZZz7gEgPnnyBBljeHJycsN3e39RAuQb4JzjNvuKV2/bZAhorUEpRW0fCPkWdoeDIyJqrXE0GqFSCvM8v+m7961JKV9KdnjvGSVHCSH77OpJ/6v/3bYtrFYrqKoK6roGxhgYY0ApRafS9ljXDosxBkop0FqD9x6apoGmafrN+dU+1R2aDUIIIYQQcr1XrZO6xMd1B0rokMmdgADQPcYREb0QouGcl0KIbvh5IYQolVJNCMEtFovAGKO2Ka8BJUC+ISFEBIDIOY+MscgYQ601aq0xTVM4ODiA+/fvw2QyAa01nXok5GvslO318z9ijNjd9qn64/j4mP3Hf/wHa9sWAABijAwRObtc1fCdShBCCNk7V1thde8zxiCEAM45aNsWEBGSJAGtNYQQYDweQ5IkoJSiddGeYYyBlBIGgwEgIjjn+pYL3YnE3eTW1SoQGpBOCCGEEHK93QMku3M/dltfSSkhSRIYjUYwGAz6w0Vkf3WJD+dcsNbauq5r51zJGMsYY9m2+iPXWlda68YY4+q63pu42G1HCZBXmM/n2LYtSClxWwGCnPMgpQxCiCCECEmSxDRN8cGDB/DgwQP213/91+zhw4fU9oGQr3FdJVWX+NhsNnB4eAinp6dwfHy8Vxd7KSWLMTLGGGdbcFkRQm2wCCF767rN1m77zy5AXlUVnJ2dQQgBqqqCw8NDWCwWfe9isj92+0orpfq5IN3Ae4AvZ3i9KtlBm3RCCCGEkFfbPVy0mwDRWsNwOITZbAbz+RwmkwkYY0AIccP3mHwfMUb03oc8z9uqqqo8z4uiKDLn3AYANpzzDBELIUQlhLB5noezszOq/nhNKAHyFbTWKIRApVT03kfGWBRCeM554JzHJEniwcEB/O3f/i28++677NGjR2w+n7PxeEwXJkK+xjZYEmFbASKlxBgjhhD2KunRSZKEWWtZjJEzxhgishgjB4Du1iVECCFkL12t/uhmQEgpIYQAbdvCxcUFZFkGWZZB27aQJAn1Kt5z3anEEAJ478F7DwBfPg+697vP7bxqhgwhhBBCyJtot+Kjs1tdG0IARAQhBEwmE3j48CEsFou+CoQOWu83RIxN04Qsy+rlclms1+uN934dQlgLIdaMsYxznocQqhBCWxQFJT9eI0qAfAVjDEopERGjEMIzxpz33gshnJTSGWPCeDwO9+/fx7fffhvefvtt0FqDlJIuTIS8wmVuALu32LWV45xHYwxOJhMMIeAeVX+w09NTBgAQQugTH4go+OWFgN+l9leUwyHkzXW1XB8A+iRId2qtrmuoqgo45zCdTvvWWGR/dXNAhsMhjMdj8N73G/SuTcPVdS8lPwghhBBCXnZ1L727hu4OmnQf01rDdDqFyWTSJz8ozrjftl1PnLW2rqoqL4piHWNcM8Y2jLFMa50zxsoYY922bfvHP/4xLJdLWlC/JvTqeYW33noL0zTtkh9Bax2klE5K2XLOnRDCK6WCMSaORiOcTCY4GAyYMYYJIajdDSFfYSf5gYyxKKWMiNi3wbrp+/dtPXz4kFlrWQiBcd53v2IAIBCRb297fU2gxAchBODlKpDurRCi35DFGPuZIM65fhNH9pcQArTWMJlM4PDwEA4PD2E4HPbJr6vDOnefG/S7gxBCCCHkS7str3YTIF2VbQgBYox9G1JjDCilQAhB66o9t+2AEhCx8d6XMcYNImbbGSBFjLGUUtacc9u2rTPGxA8//JA2Uq8JVYB8hcFggFLKyDmPIQQvpXTee6eUaqWUbjsLpBuMTk9KQr4FzjkCQGSMRcZY7JIfIQT03uMf/vAHeP/992/6bn5jxhgWY2Tee8YY47CT/ACAvR6CTgstQkhnd94D5/ylgdhCiH5WRDc3gk6q7T8hBKRpCkdHR5AkCaRpCs+fPwfvPVRVBQDQPx+EEC9t7AkhhBBCyKVXJT9CCH0FSJcM6aptyZ2CQggvpWyMMYUQIgeAXAhRcM4LpVQFAE2apu2jR4/8ZrOhWPNrRAmQrzAcDhEAEACClNIxxqwQopFSNkKIVinVKqX8NgmC24AuRQoJ+Ro7A9D79ldbfQLk/fffRwDAW37BZycnJ+y///u/uTGGCyE451xIKeVoNFJSSnN4eKhHo5HWWnPOOV0fCCF77eqw690WWFJKUEr1JfreeyjLEpIkAQAArfVL1SJkP3Rz7YbDYf9+V+HDGOtngnTPg90k2e5Gn5LphBBCCHnTIGK/Xt79WDfwvEuAIGJ/gGg0GkGapjRb+A5AxIiI0Xsf2ratrLVFjDHjnK+VUmtEzKSUhRCiCiE01tq2KApf13V48uQJzQB5jWgH+grHx8dYliUCQDTGeM65M8Y0WutaSllLKZttJYgXQoRbHqQl5NbZtr4KQogQY+ySIPjixQsAAPjd7353w/fw6yEiHB8fs8ViwbTWDC7nfYjJZCLv379v3n333cGjR4+G9+/fTwaDgRRC0DWXELLXdoPYu8PQu8RGlwQBAKjrGs7OzuDs7AxWqxXUdd0Hy8n+YIyBlBKSJIHhcAjT6RQWiwXcu3cPFosFjMfjvvJnt0Xa1SHpdIqREEIIIW+aq2ugq5Ufzjnw3oMQAsbjMdy7dw/u378P0+kUjDGUBNlziBidc64sy2qz2WSbzWZlrb1AxAut9VIptRFCFFLKOkmSxhjT1nXtP/nkE6r+eM2oAuQVnj59Cv/wD/+ASZKEtm29MaZFxEZKWWutK611I6XsWmHRE5OQb6erroqMsSiECJzzqLWOaZpi27b4+PHj2/6aYh999BEDADaZTNj5+Tnftr7iBwcH6q233kru378/mc1m4+l0OhiNRlopRQkQQsids9sSS0rZl/HneQ7OOajrGqy1LyVHyH7inEOaprBYLEBrDYPBAJbLJZyfn/c9q69Wf3R2K0MIIYQQQt4EV+fndQmQruVV27b9YaLDw0N48OABLBYLmE6n/fBzsr9CCNFa267X63y1Wl0URfECEV8AwJnWehlj3IQQKkRsYoxOCOEBIJycnFD1x2tGCZCvkGUZDofDuH0CtoyxWkpZee9LKWVljKmNMVYI4SkBQsirdQPOETF471trbeuca2OMDgA8IkYhRAwh4MHBQXz06NFevJ6Oj4/Z6ekpN8YIrbVomkYyxmSapmoymZh79+4l4/E4GQ6HRinFOa1eCCF3CGOsnwECAC+V98cYwVoLTdMAYwySJAFrLYQQburuktegG8g5Go1AStnP/LDWAmMMmqbpkyDXbfgpCUIIIYSQN8F1la+7lR/dekgpBVprmM1mcHh4CPfu3YP5fA5JkvStZcn+ijFG772rqqrMsmy92WyWxpgLrfVSa73mnBeMsdpa285mM/d///d/8fT0dC/iYfuGEiCv8LOf/QwPDg5wvV7HyWTiAaCVUtZN05Sc81JKWUopa6WUlVJ6zjll5wh5NQwhBGtta62trbVVVVW1977lnDuttQ8hRGNM/POf/wyPHj266fv7ddjJyQk7PT1lP/nJT3jbtsIYIwFAlGUplVJqMBjo8Xisx+OxNsbQkWdCyJ1z9aR/VwUCcJkAcc5B27ZgjIGmaWiY4x3AGAMhRH/rZoBYa/vZL7utznaTH7tfgxBCCCHkLrp6AKT72HUzP4QQMBgMYDgcwmKxgMViAbPZDMbjMVVN3x0xxujatq3qus7yPF8h4koptUrTdB1CKLz3dQihlVL6o6OjeHJyQhumHwClEl/hww8/RGNMfOeddzwiOgCwIYRSSpkLITKtdWaMyY0xpVKqFULQkUZCXiHGiM45l2VZ+eLFi/Xnn3++Ojs7y8uyrL33LQD4JElCCAGttV17rFs7AL2b/XF8fMyFECJJEmmMkZxzpZRSMUYVYxSIyCnQQwi5q65LZuzOBLl6o+TH3cI5B601zOdzeOutt+Dhw4dwcHAAxpg+MdY95pzzl2aCEEIIIYTcNd3hoKvJj93Kj671FQCAMQbu378P77zzDrz77rtwdHQEg8GA5n7cLcg590KIZjvsfMMY2wDAhjGWIWKllLKj0cj913/9V3z8+HGEy3gYec0oAfIKjDGYz+fx2bNnMc9zb61tvfdNjLGSUhac80IIUTDGCu99Ya2trLWNc84hYgB6whLSQ0T03vumaZrNZlOuVqsiz/PSe98gYiuE8CGEmKZp1/7qVr9+PvroI7ZarTgAiMPDQxFjVFJKHWM0AKBjjAoRBQAwRKRoDyHkTroumL07GL2bCbJbJVBVVV8hsNs+i+yfrm1DmqYwnU5hOp3CcDjsk12780AIIYQQQu66rzrs0SVCGGP9HLXdtleHh4cwHA77tTPZazHGGJxzrXOuadu2RsSSMVYwxnLOecY5zxGxBIDae99uNpswHA7jRx99dNP3/c6iFlhf4fT0FD///PP4d3/3d15KyZRSPMZYxRgLKWUupcxijFld11lRFBnnPE3TNAUAI6VkjK5ahHQQEYO1tq2qqs7zvGKMVcPhsJFStgDgOechhIBt23bJj1ubBDk+PmYAwKbTKd9sNjJJErVcLo0QQjPGNCKqGKOMMXJKgBBC7rLdAPfuqTdE7JMgMUZo2xayLOs3dYPBAIwx1Nd4j11th2WtBa01AEDf4qF7/LvH+brh6IQQQggh++5qa9ira+Tu4I8QArTWMB6P4eDgoL9Np1NKfNwRIQQMIfi6rtumaaqqqooQQo6IuVIq45xnUsrcGFMCQJOmaXt0dOQ/++wzan/1A6IEyKvhyckJPHnyJGZZFgCAHRwcNACglFJljDGPMa7Lsrz44osvhk3TqMViwReLxcF8PmdCCEEXL0JegkIIzzlvhRAWACwAWMZYK4Rw3vtorY0hhNteAdLP/litVnI8HqsQglFKGSFEAgBJjNFsq0AoskcIeSO8KhEihADvPWRZBiEEKMsSmqaBBw8egBCC+hvfMbu9rb33/XMgxvjSAPSrQQJCCCGEkH12Xfxvd/ZHCAGklJAkCSwWCzg6OoKDgwOYzWZgjLmBe0x+KDHG0DSN3Ww22WazWZVledE0zcp7vxFC5JzzwntfWmvr0Whkv/jiCw8A4ZNPPqHy+B8QJUC+xtOnTxEAwi9/+UvUWsfValWHELSUMo8xruu6Tp89e5ZUVSWdc8oYo0ajUaK1TuhUIyGXGGPIGIvb3odWKVUjYi2lbKSUVkrpYoxhPB7HFy9e3Or5HycnJ+zhw4fs8PCQL5dL6ZwzMcaUMTZAxAHnfAAAppsDAgCUCSWE3FnXnXTbrQABuAyKd62vrLUQYwStdd8KQCkFQgiqBtljuwkvpRRIKfuTjlcrQHafI5QEIYQQQshdct1hjxACOOeAcw5KKZjNZnDv3j1YLBaglAKlFFV/3CEhhGitbTebTbZarS42m805Ii4Rcc05z2KMBWOsTNO0EUI42CY/ttUftDD+gVAC5KshAODTp0/Zz372Mzw+Po5CCJvneR1jLEIIG+dcmud5aq01WuvRw4cPJ4g4A3rSEvISznnknDullGWMWc55s33bMsb8eDwO3nt8/PjxrX/tzOdz9uLFC5GmqQwhaABIGWMDzvmAMTaIMSaIqACAxxgpokcIudOuBrG7GSAAX558896Dcw5CCCCEgDRN+wTIeDwGrTUlQPacEAKMMTAajaBtW6iqCpxzL7XDAvjyhCQlPwghhBByl+weCrpu+Hm3HkrTFMbjMUwmkxu+x+QHEhDR1nWdl2W5zrJsqZRaa60zrXURY6wAoPmf//mfFgDCkydP4gcffABAceQfFCVAvhk8OTlBRGT/9m//FowxrZSyqqoq55wnbdsmQoiBlPJAKdUAQLitp9cJuSHIGItCCMc5t1LKmjHWKKUaIUSrlHJKqTCbzSLc8ov+8fExK8uSc85FWZaKMZYg4gARh4g4AoABIiYxRk0VIISQN8XuqbVuwwcAwDkHROwHYyMi5HkOf/7zn6EoCiiKAt5++22YTqfUDmuPMcbAGAOz2QwAANI0heVyCavVqh96L6Xsnw+UBCGEEELIXdOta2KM/fqmS4A450BKCc65l9bK5O7pYl9KqVIIkXHO11LKjRAiF0KUQojGe+9gm/yg+PGPgxIg3wJjDP/1X/81SCmdMab23hcAYDjnKed8xDnPt0PS7fbJLDjn3TB0CoKSNw1uf/ljuOQAwAohaiFEzRirtda11toiotNaB+89Aly+1m74vr8KOzo6YqvViidJIgBAIaKJMQ6dcyNEHIYQhoiYhBB0jFHQEHRCyJtiN7AN8GVSpAt6SykhhABVVUFVVdA0DXjvYTqdwmAwuKm7TV4Dznk/0FNr3Q+7t9ZCCAGapnnpNCTA9cmPq88hQgghhJB9sFv90ekqP7rWsFJKEEL07UDJ3YE7QgguxtgwxgopZaaUWnPOM2NMzjmv0jS14/HY//KXv6Tkx4+IEiDf0nw+jwDgpZQ2xliFEDTnPEXEUYxxXVXVZrPZZDHGNE1T0FprKaVgdHUjb5jthT9677211lZVVTvnKgAopZQFY6wUQlRa6xoRW2tt8N7f+gqQTz75hB8cHEjvvWKMaQAYhBBGIYSx9368TYakIQS9HYJOr31CyBth91Q/wMszQbrkR4wRnHNQVVU/C6SbC0L2W7epT9MUGGN94qNriea9/4sEyNXKIVouE0IIIWQfXLduudr2qqsEkVKC1hpGoxFMp1NI0xSEEDd0z8kPARGj9963beuapimbpskQcc0YWyml1mmaro0x+XA4LBlj7XK5pM5BPzJKgHxLp6eneHBwEN977z2X57n13tcAUMYY8yzL1p9//vlFXdeT2Wwm5/N5PDg4mHDOE7q4kTdNjBG99z7P86YoiqKqqqxpmsxamwNAAQAlANTWWqu1bquqClLKWzv8HADg448/5mVZ8rquBSKqtm1NjDENIYzath1774cxxkEIIQkhKESkChBCyBvnaln/7iBIznk/LJtOv9093ePZtcNCREj1PKL0AAAgAElEQVTTFC4uLiDLMqjrGpxzfUu0q8+B7rlCyRBCCCGE3FZX1ynXzfzw3oP3HpRSkCQJHBwc9LfZbAbGmBv8DsjrFkIITdM0WZaVZVkuq6q6yPN85b3fcM4z51ypta6dc1Zr7e7du0env35klAD5lj788EP89a9/HUMIPoTQxhgbRKybpikQcVPX9fl6vR4dHh5qRORaa8M5lwDAGGNsOwCSdnTkzkPE6JzzRVE06/W6KIpiE0LIEDEXQhRKqVIpVQFAwzl3dV3f6uoPRGS/+93vWNM0wnsvQwiqbdsEAAbe+1EIYcQYG0sph1LKhHOuAYBmgBBC3ji7J/x3dQkQIQQIIfo2Sd0m0TkHnPM+SUL2l1IKRqMRKKXAGNNXgHjv+1YQX4eSIIQQQgi5ba5bn+zO/thtewVwWSE7HA7hwYMHcHR0BPP5HJIkAa31Tdx98hrh5YOM2xkvrizLerVabbIsW+Z5vowxrkIIGwDIhRBFjLH23rfW2vD+++9TAuRHRgmQb2l7YQv//u//zkejUVuWpRVCVN77smmaTVVVq6qqRgBgjDE6SZIEANhgMEiSJJGMMWqHRd4I2xZYwXtfN01TlGWZcc4zKWUOAAXnvOSc1957yzl3xpjw2Wef3doEyNOnT/loNBKccxFCkCEE7ZxLYowDRBxJKcda65FSajSbzQaj0cgopQTnnF7vhJA3yqvaGnHOIcbY90BmjIH3HoqigM1mA0IISJIEjDEgJS1R95kQAowxoLXuH+e6rgHg8vnRtm3fFqLri02VIIQQQgi5za6r/AC4HHS+m/wAuFwLaa1hOp3CYrHob+PxuD/wQ/ZbjDE652LbtqGqqnq9Xhfry9O/67qulwCwYYxlWuuCMVYBQDMYDNo8z/3Tp09vbezrrqLd5beHAABpmoY///nPjjFmhRCNc66MMWYhhJW1dpDnuT47O5OIKIuiiIvFYrxYLIZJknDa1JM3AWMscs49Y6wWQmRCiDVjbCOE2CilMs554ZyrtdaNlNKt1+t4enp6K38JdNUfZ2dnvGkaGULQ3nuDiIlzbsA5HyVJMp7P59PFYjE9OjoaHx4epoPBQAkh7sTK5mpLG0II+Sa6AegAX1aASCn74Le1Fp4/fw7OOajrGg4PD2E6nVICZM91bc4ALtthTadTiDFCkiSQJAksl0uo6xratu0DAF1brN2vAUCVIIQQQgi5ebtDzq9rf9UlQbz3oLWGwWAA8/kc5vM5HBwc9JUfSqmb+hbIa9a2bSzL0q5WqybP8yzP81VVVStr7RIRV4yxtVJqwxjL27atpJTNF1984R4+fBg++eQTCq78yGh3+R0wxvDk5CQeHx/7Z8+eOSllkyRJhYiF934DAKm11pydnamyLHVZlgwR2WAw0FprBZdtcQi5i7ZVgJcFIIyxVilVaa1zY8xmmwDJhRAlAFRCiBoR2yRJXJqm4cMPP8STk5Mb/hauxc7OzjgACOec5JwrRNTbWR8pIg6VUqP5fD76q7/6q/Hh4eFwMpkkxhgppdz7qA0lPggh38XVE/0AX1aBdEmQpmngxYsXUNc1WGtBKQWDweCm7jL5ASilYDgcgpQSjDGglAJrLTjnoG3b/vNijH8RUKDTkYQQQgi5adfNtus+3iU/dt9KKWE8HsODBw9gsVjAfD6HNE2p7dUd470PRVG0z58/LzebTVaW5ZpzvuKcr5VSGwDIGGMFbGNfZVm2z549c//v//2/SBUgPz7aVXxHJycn8fT0ND548MBZa1spZaO1LrXWGed87b2/KIpieX5+vtxsNpu6rqsQggMA6vNG7ixExBijb9vWWmtLa20WY1wDwFpKuZZSZlLKHBErznkTY2yFEC7LsvD48eN4GwegIyJ7+vQpOzo64nCZvFQxRh1CMF0CxHufMsbSJEmS6XSazGYzPRgMlFKKUwssQsib6upmsbvtlv2HEKCqKiiKAvI8B2stxEhLpbuka4c1Go1gOp3CbDaD2WwGk8kEhsNhHwzoTk4CfFktRNUfhBBCCLktdpMfAPAXba+6Qx/T6fSloeeTyQSMMX11LLkbQgixbds2z/NqvV7neZ6v27ZdA8BaKbVOkiTXWlda60YI0U4mE/fFF1+Ep0+f3ur5t3cVVYB8PxEAwng8dm3bWkSspJQZAChElE3TaM556r0fxBgnjDEP9CQnd9i2B6Kr67qs63rVNM25tfYCAM6llEvO+YYxVjLGqtFo1EgpW865/9Of/hSPj49v7Wvj6OiIFUXBAUCEEGSMUTPGTIzRhBAM59zEGDUAaKWUlFIKpRQlmAkhb7Sr1WNdMHt3GHoIoW8X0A3IpgTI3dK1w+pmvEwmEzg8PAQhBCilIM9zqKoKnHN/kfTYfUvViIQQQgi5Kd1aZHfgOSJCCKFve9Wtc+bzORwdHcFsNoM0Tant1R3FGAsA4GKMVQghb9s2S5JkzTlfCyEyKWXJGKsHg4H13rskScLJyQltdG4IJUC+hw8//BB//etfY5ZlnjHWJklSCyEkY0x476UQwnDOR1rrqTGm5pwHoAQIucNijKFtW5vn+Wa9Xp9XVfVcCPGcc94lQDLGWLl9PbTD4dBfXFzEx48f3+pfAuPxmAEAX61WkjGmEFEzxgxjLNlWgRjvvfbeyxgjR0Q6rkoIeeNd3SheTYB0LQK6llhCCGp5dMdJKWE4HML9+/f7gfcxRrDWQtM0AADXVnxQ8oMQQgghN+HqTLLuoM7u3A/nHBhjYDwew1tvvdW3vRoMBpT8uMO2c2+dEKIWQhRSyg1jbM05X0spM855BQC2KAofQojOOVrQ3iBKgHwPjDH4+OOPo9Y65HneCiG4lJLHGJnWWnjvNQCMGGOjtm0nZVkutdYCEaOUUnHOBWOMauDIXrvsehWj995ba6uqqrI8z5dZlp1VVfU8SZIXg8HgTGu9EkJknPMSEW1RFO6zzz4LABCPj4/xNra/AgD46KOP2PHxMQMAoZSSQghtjNHW2mQwGKSDwWAgpRwtFovhZDIxSilBba8IIeTS1WD27un+rhVWl/iIMUJZlrDZbEBKCVpr0FrTQPQ7RAgBjDEYjUb988BaCyGEPqjQJcs6XdKMkiCEEEII+bFcPcQDAH8x6wPgsu2V1hpmsxksFgs4PDyEg4MDGA6HfQUsuTNwG/uKzrlYlmVd13WJiDljLAOADed8tU2CZFLKChFtmqaurutwdnZGi9kbRDvK7wdPT0/x4cOHwRjjtdYtAHBEZDFGKaVMEHEVYxzUdT1cr9cDxhgfDoc4Go1GSqlE0NWQ7Lmu7VVVVU1d13me55uyLFfW2gvv/YX3fhljXHHON1rrgjFWO+dazrk7OzuLp6en8YMPPrjVvwhGoxErikK0bSsBQDHGjFIqGY/H6WAwGA2Hw/HBwcHo4OAg1VpLSoAQQsiXdis/rrY36hIgiAjWWliv1yCEAO89zGYzGI/HfdCc7L/ddljdqUlrbV8NVFUVNE0Dzrn+8wGoAoQQQgghP57ddcfVgeddu9augjlNUxgOh33iYzqdwmAwAGPMTd198gNBRPDex6qqXJ7nbZ7nRZ7nuXMuB4BsO/h8I4TIAKAAgMYY0woh/Hg8Dp988gktaG8QBd+/p9/+9rfw6aefQpqmXRYYGWNoreWIKKSUAhGF955VVQUhBM4YE0mSJFJKJYSgJBTZa9573zSNXS6X+XK5XGdZdtE0zVmM8YUQ4kxrfSalXKZpuooxFk3TNFJKe3Z25quq8v/yL/9yq38J/PM//zNfrVaCc24452nbtiNr7dQYM5vP50dvv/32W3/913/9Vw8ePFgcHBwMh8PhnRl+3jQNlGUJWZZB0zTQtu21n0eBSULIV9lNfOxWfwC8vKn03kPTNGCtBWtt30s5SRK6ztxRUsr+5KRSCrz3YK19KQGy+7zpPkYIIYQQ8kPbXYPstrzq5tZprWE+n8Nbb70FDx48gMPDQxgOh6CUoraudxAiorXWbzab5tmzZ+X5+flytVqd13X9IsZ4xhh7obU+M8asjTG5EKJmjLXz+dydn5/Hf/qnf4offfTRTX8bbywKvn9PjDE8OTlBAIgHBwf+nXfewe0gTymE0N771HtviqJQRVFIzrmSUsokSRJEZIgIQgjJt276+yHkm4gxYowxhhCitbapqqoqiiIry3JVVdWSMbbknK+klGul1EYplQkhSqVUo7W2WuvdDPitToAAALRty40xwnsvQwiac64ZY0mSJOl0Ok0Xi0U6Go0SrbWWUt6J5AchhLxOV1sYXa0C6TaTzjlAROCcQ9M04L1/qWqE3B2c834mSBdUWK/XfSus6yqGAKgahBBCCCE/jG6NcXXNsZv8ALg8wCGl7AeeHx4ewnw+h+FwCFJKSn7cYSGE0LatLcsyz7JsU9f1GgDWiLjRWmdCiBwRyxhj3bZtOx6P/WaziY8fP463te37m4ISIK/ByclJPDk5gQcPHuDnn38eAQDm83lVlqVs21Y750RVVTyEwC4LP6QUQhjnHDjn2Gg0SrXWmhIgZF/EGGPbtr6u67a6lFVVtWzb9sJ7fy6lvBBCLLXWK2PMOk3TTEpZTqfTZj6ftwDgHz16FH7xi1/c6uHnAACnp6fs3XffZXVdixCC4pxr732ilEo454nWOhmNRno4HFJFFyGEfIWrQ9EBoB+GDnC5uXTO9RUgXTKE3E3dDBgpJYQQoGmavk92COGl4MF1lSAAlAwhhBBCyOuxe+ji6vqia3+12/ZqNBrBbDaDo6MjmM/nMB6PQWt9E3ed/HgQEUOMsWnbNnfOrbz3SynlSgixFkJslFJ5kiTleDyu27ZtP/300wAA8f3336dF6w2jYN1rcnJyEhGRffTRR/jw4UMAAG6MqbXWeV3XknMunXPCWpssl0tT13VSFAU7Ojrqij+EpCmfZE+EEGJd1+16va7Kssyqqlo751aMsZUxZqWUWmmtV0qpTYyxaNu2unfvXl2Wpfviiy/C8fFxhD2o/Ojkec7SNBVCCOmc04wxAwAGEU2MUcYYOSLS8WRCCPkWdhMiXSAc4MtTdTT7483SBRZCCOC9758Tr0p+EEIIIYS8LtclP3aHn4cQAABAaw3T6RQePnwI8/m8n/lB433fDJzzoJSyaZrmdV1vYowbKeVGKbVhjBUAUG02m4ZzbsfjcQCA+OTJE6r+uAUo4P4adU/ojz/+OJZl6WezmXXOVUIIWVWVZIyJGGNSlqWuqkojIlNKicFgwDnnyBhDaodFbqsYY0TEuE1+2KqqyqIosqqqVnVdLxljF0KIc6XUhVJq2bW+AoDSGNNUVeWeP3/uP/3003h8fLw3vwAePnzIAECEEGQIQYUQTIzRhBDSEIJBRIWI9HolhJBv4GoQeze43QW8uw1k27ZQFAUkSQJa676lAAXC7x7OOQghwBgDaZpCXdcvBR26ZfHV4ESXRKM2aYQQQgj5Pq62awV4eb3RrUW7tleLxQJmsxmkaUozP+427OJg3vvWOVciYiaEWCulVsaYlRBiI4TIlVJFCKEej8cWAPxvfvOb+OGHH+K+xL7uOkqAvH74q1/9Kv72t7/1RVG02wHo3TB03jSNbttWtm0rOec8SRKZpqmAyxcVDgaDVGutAICunuRW6dpeWWvbsiyrsiw3dV2v6rpeOufOtdZn2wTIuZRyJaXcDIfD3FpbI6J99OiRe/ToUfzFL36xF3M/tpi1lkspOSLKEILeJkDSEELivU9CCAoRqQKEEEK+pd1N5W4rLMYYhBCgKAowxgDnHMbjMQwGA9BaU6D7DuoCC8PhEGazGYQQoK5raNu2rwy5WgnSJT6oDRYhhBBCvo+rbVqvrjG6QxqDwQDm8zkcHBzAbDaD0WhEba/uOERE73303tuqqqq6rrOmadYAcKGUuogxLrezbzOlVMU5t3meu3/8x3/0AAAnJyc3/B2QDtVo/UDeeecdmM/nEGOEoigAEUFKGbcXUWSMIec8xhixqqronIvee3Y5Q1kqaodFbhtrrSvLsrm4uMjX6/Uqz/Nz59w5ALyQUj6XUj7jnL+QUp4rpZaMsbW1thiNRpWUsp3NZn6b+d6HSAUDAIaI7D//8z+1cy5BxAkizpxzByGEBef8cDgcHs7n84P5fD4zxiTijtW9Nk0DZVlClmXQNA20bXvt51EwkhDyXVy9duxWd3QzIaqqgrZtgTEGxhjQWtMJuzsIEUEIAUqp/nH23oNzrk+CdEvjV/3OuTo0nRBCCCHk67xq/bDb9ipJElgsFvDw4UO4f/8+HBwcwHA4pMqPNwAiRueczfO8uLi4uFgul883m83/1zTNn2OMX0gpXwghLqSUGSIWMcbmj3/8o//Nb35z6+fdvmkoyP4DOTk5wY8//jiMRiPXti2v65oLIRjnXF3OQBecMcaqquLW2m6QDo5GIy6lRESMcBmE5YwxLoTo/j7bfpyQHxoiIsZLwVpblWVZZFm2KYpi1bbtuZTyvKv64JyfAcCSc74KIWRCiEIpVWdZ5pxz4Z133tmb5MfJyQkDAP706VMOAEoppZumMQCQKqWGSqnxYDCYjEajkVIqYYxJoNclIYR8K7sn97tNZ7cJ7YLfTdOA974PjDPGIEkSmhFyx3SP5Xg87ud+tG0Lzrm+AqRzXdXH7vOAkiCEEEII+Tq7FR8A8BdrjRhjP5OMc95Xqc7nc2p7dcdt42AYY4zOOVdVVZ3neb5er5d5np+3bXsGABcAsJRSboQQufe+SpLEPnr0yJ+dnVHy4xaiBMgPB3/1q1/Fjz/+2Dvn2HQ6Zd57YIwJROSMMdY0DXPOMeccxhgRAGA+nwvGWLDWuhijhMvgq0zTVBljJOf8Tp0wJ7fX9pd+cM65tm1tWZZ5VVWbPM9XZVleeO/PRqPRmVLqQmt9zjm/kFKuGGMbxlhZVVWdJImVUrqf//znAfYk+QEA7PPPPxd///d/z5umkUopXRRFAgApY2xgjBmlaTodj8ez+Xw+SdN0IISQjKIthBDyre0Gq3fbDsQYoWkaALjckBpjQCkFMcZ+2CRjjAZO3hFdcEFKCVJKQERomgacc8AYg6ZpIIQAMca/GE56Xc9uQgghhJCvcl3lx+46NIQA3vt+ram1htFoRG2v3gwYQgh1Xfu6rpuqqsr1ep1tNptlURQXIYRlkiRLpdRaa50xxkpjTD2ZTNqLi4vw5MkTSoDcQpQA+WHh6ekpAkB89913vRCibZqm2SYxmNaahRC4UgoQMTZN458/f+43m00upZw651Kl1CBN08HR0dFgPp8zKaWgOCv5kaD33td1XWZZlm02m3VRFGvn3JIxttRan20rQJaMsSVjbIOIRQihBoDGOddeXFz4NE3j8fHxvkQm2MnJCQcAUde1GgwGKoSQxhiH1tpRkiST0Wg0e/DgweLw8PBoMpksxuPx2BijttVZhBBCvoXrTu53NyEExBihbVs4Pz+Htm0hz/O+/cDuwHRyd3DOIU1TWCwWIKWEwWAAq9UKlstl3w6ra5d2dRg6VYIQQggh5Ku8KukBcHnopqv86KqRQwj9290qEXJ3xRixbVu/Xq/r5XJZlGW5qqpqaa1dMcZW3cwPRCxjjLXW2g4Gg3YymYSf/vSn9CS5pSgB8gPrWmE9e/aMzWYz0FpzAMAYY2SMRSEEMsZ8CMHVdd2cnZ3VnPM5Ik5DCGNjzHQymUy11sEYg0opEEIIxhindljkNelaXSEixu2MmoiIwTlXVlW12Ww255vN5qKqqlUIYSWEWAohzre9DldKqQ3nfMM5L621ddu21jnnfv/73wcAiB988ME+JEDYkydP2MXFhUjTVGmtdVVVqfd+3LbtxHs/iTFOlFKz+Xw+Pzw8PBiNRjNjTCqllIwxqn8lhJBv6brT+91QdCFE3w4ryzKo6xqcczAYDGA2m/XtB8jd0g0anc1mYIzpW59ZayHG2LfF2g1gXK0kIoQQQgjZtbvejDG+MgkihOjXod2BnG0cjlpevSEQEdu29XmeV+fn55s8z5fOuYtt6/cLrfVKSplJKQvnXC2ltADgLi4uwk9/+lPczr4ltwwlQH54fSus0WgERVFYAEBrbQwhxCRJ0DkXGGPOWtvUdd3EGEvvfYGIszRNXYwxzGazOBgMUGuNxhgjpVSMMUmbPPJ9ISKEEKL33jvnPCJ6zrkHANc0Td627UVRFGdVVb1wzi055+vtBX+plFpqrTeMsRwASillLYSw8/nc/elPf/IAEE9OTvYiA35ycsI+//xzvlgsxLbdnHHODWKMoxjjpG3bSZqmE8752BgzHg6Ho9FoNBBCUP0rubV2T0d3XjE+uPsb3+7rv/of/lZf58551ZDm1/TlEeDLn/EerwOuS37sBra7tkjdQHRrLUgp+0QItT26mxhjfSssrTUwxsA5B1VVQYwR6rqGtm0hhNBXg1wXkNhNjhBCCCHkzbXbMnP3wETXWrNLiHDOQWvdH7Bp2xaEEDCZTPoZdBSDu/sQEUMIoW3bOs/zfLPZrBFxORqNlsPhcKWU2kgpCyFEJaVsrLXtdDr1x8fH+9L6/Y1ECZAfBz558iQ+ffrUP3v2DN55553Ytq3nnAchRAAAJ4RoAKBCxGqbAClDCE2SJA4AbJZljRCiCSG00+l0Mh6Ph0IIDgDU+4F8LzFG9N77sizrsixr733NOW+klFUIIbPWLqWU50mSnAshVkqptRBiLaVcCSHWMcbCGFMiokVEZ4xxFxcX4fHjx/GDDz7Yi+RH56233mJpmgrvvU6SJHHOjRBx4r2fee9nTdNMrbUj51wSYxSISKsfcmtd7Y3flQwi4mUgvl+8f83TeDd4eGXBz+D6FR4y1v+9N3KTsPP9v/Th7/Cl+scLvvxZc8YAu8cWERD29+d8NQmyG7TuTt/FGPtBk93brgUSudsYY301SIwR0jSF5XIJy+USvPcQQgApL7cz3XPiujZYlAQhhBBC3lzXrRmvVoRIKcEYA4vFAiaTCRhj+sRIkiQwn88hSRKqAnkDMMZQCOGllI0xJhdCbBhjK2PMhVJqKaXcaK2LGGMzGAzaxWLh//SnP8Xj42Oq/rjFKAHyI9m+COKTJ0/8crkMx8fHvmmaMBwOPQA4zrkVQjTe+yaE0L11UkoXY2zzPG8QsUFEJ6UMxhjYts+SsI2pbIOxbLv5Y5xzth3MTBECchXi5W/8uM1sN2VZFpvNJrfW5pzzQimVA8AGAJZCiOVgMLhAxI0QYiOl3HDON1LKzDlXK6WaJElclmXhpz/9aVf2t1fJj+PjY3Z6espjjDJJEm2tTQFghIgzIcTcGDM3xsw45xMASICun+SW2734MwBgO4kQ6IPqDBjg9VUEuxUG2yD7S8H2yw+8/G8ydvnn132dV9iX4P1LQfpv8Pldsukv/s7VYOx1P56df+ClLRbiS8mVPpGF+OXjsQc/y6t2A9S7VUvdBnP3ZF73uc45cM6BEIJaEtxh3UnM0WgEUsr+RGbTNOC97z+PBqMTQggh5JvYrTbuZn50ByqUUjCbzeDo6Agmk0m//uySI8YYWnPeXdgJIfgYo2WMVUqp3BiziTGulFIrrfXaGJNJKSvvfd/66vHjx5GSH7cbBfB+XPj06dPw9OlTAAD4+OOPw9HRUUjT1Gut27IsbdM0NoRgEbGu69o652wIoWqaJvPe54yxejAYtMaYNsY44pzrGKOIMQoA4DFGIYQQSilhjJFCCEHDmclVlyM/LnMf29ZrRVEUmzzP19baNQBsjDHrnWqPtRBizTnPpJQ557xgjOXW2hIA7HvvvdcCQNzeYB8v/KvVig+HQ2GMkWVZGgAYeO8nQoiDJEkOjTFH4/H46ODgYJ4kyYBzLtk+RG3Jm6UbIt39d4yX1QLbhMeXyY/L//UB9X6g305ZOMBLSY/ucxEAIOJO16wvg+59tcJLiZK/PN3f393u/7p/4xZXDF89TXBte53u+4sRYPs4dD+P/s+7TddXpVG6L7n7M+7fRcCdU+5fBnsv/wLu/lt75Oqp/d2Pc877U/6ICHVdw3q9Bs45jMfjfhYIDUS/exhjoJTqAw+MMfDeQ9M0AABQVVXfDq07vbn7dwGoBRYhhBBCLu2uN7v2VyEE8N73VcZd5enBwcFf/D3a/t9dMUaMMQbnnGvbtmyaJo8xbjjnK6XUkjG2NMYstdZrIUTBOa93W1/tYwzsTUMJkBv05MmT+Ic//CG0betijGzn9GN0znkppQ8htDHGEgCyGGNurS2Loig456s8zyeImIYQTAhBxxgVIipjTDL6/9k7l95IrjNNv9+5RETebySrSi0DgiH0gmr0Rt40MEC7gdnMYLbln9B/Q9TfsbZezWJgr7rRDcOrrsEYDaNhqCWLLDKZ17icyzeLiBMMZrFKkq0Wi+R5gGRkRkZGXhmX7z3v+w2H2XQ67WVZRiJK1JEDmNk756r9fr/e7/fr3W53XZbltff+mpmvhRDXAJbMvPLer4UQayHEOkmSnZRyx8x5r9fLx+NxtVqtLB62+EFnZ2dUlqVwzilrbUJEaVVVfe/9OE3T2XA4PHr+/Pmzo6Ojk/l8vphOp8M0TTUOBmdHIvdGEDi67oCO6NEKHxxuM8C+MQzQG44Nxo2Q0ugTqPUS7ggjd/eiCLFM3fXdXD2IxeLbDpAffOPxQxU+D4ScIDrQXct0XBo3nyDQdcy038ehIHT4WbUnW43wEW40b42pjhsLrhum2tPju6/jAXJXRrMQAt57VFXVxh/t93ssFgucnJy0cVmRx0n4DYSiBDMjSRKsVitcX1+jKIp2FGf3d+D9m2ZUvuN/LxKJRCKRyOOlu+8Pgya67g9jDLTWcM4BuO1EjjwNmNlba6vtdrvdbDarzWZzsdlsLo0xSyHEtRBi5ZzbSCl3RJRPJpNqs9nY8/Nzf3p6ynifR/JFAEQB5F5pTvDdb3/7W1RVhe12y8459t5bKaUBUAkhSqXUlplHRLQxxmxXq9V6t9sthRAj5z60rWQAACAASURBVNzQOTfw3mfW2oyZ0/F4PDDGDNM0ZSllJoQIhek3XsO7ehjcUZj50c8Wv8sJ6vveh+FtgsAPOSLx256jez8RcZ16Ve3zPF+u1+vLzWZzaa1dAmhdH02/jzUzb5Mk2RLRHkA+Go1yY0yltS632639+OOPHR6u+IGzszP6+7//e/H73/9eCiFUnudJURQ9a+2AmcdSymmWZYvj4+Oj58+fH02n01mWZYnWWkd3VeS9gLmNt2qdHp2pDMX4dl4tgNRCCN04FDrF9rAugG4im5qCv29ilm45Dby/dcTXnmQcRGYFl0dX8AgyQqf0//3e/rd8Nj8IraBxs9rwORGo49QAWmPNzcNA1IaN3QhUbYzYW146uPO518/BADw8gKYHiBAA1YIHN+u7+SboQRd6uyKIEKKNK7DWYrVaYb/fI8/zti+EUqrtDRJPWB8nRIQkSTAajZAkCZIkgVIKVVXBe4+yLN8Qz4DbkViHzqlIJBKJRCKPj8P9fDcasyt+hH5i3eXi8cGTgptzDDbG2KIoytVqtVkul1fX19evrbWX1tolEa2klGsp5cZ7v0/TtMiyzIxGI/fpp5/G6KsHQhRA7hcmIvzyl7/0P/3pT+0333zDg8HAHx8f2+VyabMsq5IkKXe7XU5EORHtq6rKrbU7Iloz88h7P3TODZm575zree973vthmqa7PM9zpVSPmZPm+ajbJyQIB8zc3u7O7/DGHuAty33rfe9a560Ppnn8UxFA7lqGiPgdIsktQaO7znC7mYYmTAyAGzGMrbWlMWab5/nFfr9/nef5awDXRLQiopUQ4lopdd3EXe2NMflwOMyFENV+v696vZ7Zbrf2o48+Cu6PByl+MDN98cUXdHFxIQaDgVqtVtp7nwkhesw8cM6NnHMTIpqkaToeDAbD4XDYF0LIpsfOfb+FyFPmoLk5AJD3IACCGeS5nrIHeb4ligjcdoiIUODvFg3b4v2N4wCdmn13y3srIqtxPoRQq1tZ/N3/mUMBgNE+pl3nd4HuFhP4+wgp71j0UKpp31fzHoOQFBwyITyMcPP5UbsG3Lp2F77bC6Nt49U8EzUyihC1+CEkPBFICHj2YKqbQHs038+D2yrf0P0tBvcHEcE5h6qqUBQFmBlpmqLf77fRSFmWIUmS6AZ5hIQM7uAECbEVeZ63BYtQ0AiC2eFxVIzDikQikUjk8dK6tO/oBRaOC4LrwzkH7z2EEOj3+xiNRhgOh2j67d7TO4j8mHjv2VrLxhiX53mx3W536/X6erVaXW42mwsAl1LKpRBi5b3fSin3AHLnXPVP//RPDoD/9NNP48HlAyEKIPcP/+IXv/AvX77EJ598wqenp/7i4sIdHx9bANV6vTb9fr8siqIQQuTe+721duu9HwIYOOcGzDx0zvWZOWPmXlmWg+1227++vh5WVZVqrRNmFgAEMwtmDpVbEQSRcCEi8t5TQxAX2utBJGloBZQwoxl1+cb87yKsdEblBaHmW10rzahQOlzHX8q3iSrvKvYf7miJiEMEw6FYcbA+Pnwc2rrirbs4KCNExETEQojuPN88jonICyEcEbkwJSLHzIVzblcUxZW1dum9XxLROqjaSqk1gDWAvRAi11qXZVlWJycn5ujoyAJw//Zv/+Y/+ugjjxuR5UHy05/+VHz99dfKWpsIIbIkSXpFUQyZeeScGzciyAhAT0qZKKUkET3J4cXdA8m7DiojPx7ciBjNjVrUYK4FEO8hvAc5B+Hq2+QcJDPgfb2sb0QQ1LFYgqgWQeoV1tvSpq8EURAzbsr3YQvJndfT/ia6hfeOC6S9jdv9L/jWFb497ztA4i7x43Chb1nJHU94u09HJ7qq8/5ah0f3zmYGhX4crVukMwqts9bb7/9mHncknHqjTmDRuCEEAVICUsNLAZYSLAQceXhBIBFEEHrzeR4Ad21bghNECNEWuouiwNXVFbz32O12ODo6wsnJCYgonrg+Urrfba/Xw3Q6bV1Ay+US6/UaRVGgqqrWCRSmcdBCJBKJRCKPlzvqMO28MGgiTEPslVIKWZZhPp9jPp9jsVhgMplAa30fbyHyI+Oc47Is7Wq1Ktbr9Waz2Sz3+/3roijOvffnRPSaiK6UUtdCiI1zLi/Lsvryyy8tAPfy5cvo/nhARAHk/YC/+OIL/8UXX+Ds7Myfnp660WgkNpuNHY/HdrfbVVJK45yrkiQphRCFc26PuiDbt9b2iagHIGPmlJl7+/0+Oz8/72mtE6WUZmYJQHanRBTEkDdEkSbah5p5BIC896IjcFCz3KFb49b8rmDSXe5wfjg57QgP7Vnq25Y9XK7zGu7+kL+DU+SO9b9z8eYxt2YeOjcOb4cbYRKWCdNmlCt3HtfWGMN9uBE4GIBvlg8bX9/M80TkpJRWCGEAWCGEkVIaZi6IaG+MWTPzJkmSNRFthRC7JEm2SqltkiRbACUzl1prs1qt7PX1tTs6OnIA/M9//vMHLXwAwC9+8QvxP//n/5TPnj1TeZ4n1trMOdcXQgyEECMhxAjACECfmZPm/ycSuXe6GzMKAoj3EM6BrIOwDsJaCGcBY+p53kOwh/C1UCJQO0YECQjUDW2IDrajjaMgCCAMbmv8fLi9bR0ioehPOHRhMFoN5OAN3RYxvo/74/BB1PTEOOSdjpB3CSCEN+Qa6ggdXTnjJs6rI57cYX65cYp0nDTcFT8A1whHvnHqeCKwFLXLQ0lAKUA7CK3BGvCCASlAJOA8WqHEe9+6hR5KT5BwwtrZ97ej+ZRSt7Kb1+s1drtdG4c1GAyQpuk9v4PIj4HWGsPh8FaD9KqqbjVFP/wtBaKIH4lEIpHI46E7SC/c7l7vxlx1nSBSSgwGAzx//hwnJyeYzWbo9XpIkuTNJ4k8Orz3vigKe319nV9cXGw2m82SmS+996+VUq+llJdSymshxIaI9pvNpkzT1Lx69cqenZ09tDFmT54ogLw/MAA0/0TEzP6LL77wAPyHH37ovvzySw/AOueMlLJUSu2dc1lVVRkR9ZRSKRElxpjUe58WRZFYa1Mi0lJK5b1XQgjJzAqAEkJIABKAJCLhvZdCCGJm0agc1IxyJzR1seb+VhQJ04MIrTaNheoKPjVFCwIA7317X9ghhSsdNwrCtCOa3Kr3tVe6dpQDoeWQt7hQ7lruuyzTbujuaLDJh9e7LpAwr1E3bgkg6Lg7cCNwhHlhHcz1F+WBOtaKmX1wfgghHADHzF4IYYnISilLZjZSykoIUQkhCiIqhBA7APskSXZKqb21NldK5UqpfDKZ7IuiML1ez+R57gC43/3ud/7jjz9+NCr3J598QlJK6ZxLiCgjor73fpgkyShN05EQYjKdTsez2WyYZVkqpRQHLqhI5F4IxTsRYqw8144P6yCMgTAGVFUQlQGZ5mJtLYI0AohsHi+JagGkcYGEmn4tJDQ5uE29P0RgcRt3hXaLfNgLIzRSDw6QIIwcvo9m8Zt1HPDWjc1d/4Z3CRmda9+64Tp8fV0BpBU8Ou+18wFQ5xluvQ/u+GfC53jwPoLUHRRsRh1j5pvb4ZTNC1E7P5QC6QSUMeAY7Bki0SBC7QBpYrBc4+7x4Tt4QH0Puq8ziB/B+RGaVIbRe7vdDkmSYLvdtv0gIo+fEIelVH06Y4xphTBu+sUEoewuF8ihCPKQ/j8ikUgkEonU3JVQEK6HY4LgIlZKtfdZa9Hr9TCZTDCfzzGbzTCZTCCEiE7iJ4L3npnZlGWZ7/f7zXq9Xmmtr6SUl0mSXCqlrqWUa631rqqqot/vm3/6p39yUfx4mEQB5P2EmxMwx8z861//2u92O/7ggw/sfr83xpgyTVMNQGutE6114r3XxphESqmFENp7r8uy1EIIxcyaiJSUUhKRIqJWEEEjgjQj2wUA6b0XUkoK7pBGrLglinRFkE5M1hsCSHO9nReaRncqyIdukVZM6RSabzlEDmO2Dk5mbzlHDj/Y71K5/i4FbiHE2zZ2N2kmnZgqANzsRLnZCbOUshU0qHF8NKMQWsGj/ng53NcKIkHsoNrl0To+mNkzs2uEDwfAMrO11pZEVAGo0Lg6hBClECIXQhRpmhbe+3IwGJQAKiKqpJTlRx99ZF+9euXPz8/9b37zG392dvaoqkqnp6cCgMrzPAWQEVGfmYdpmo76/f5kMplMZ7PZZDabjcbjcaq1VrE4EnlfaDeiTfRV6/qoDERZQpQlKFyqCmQMhHOQnkGuFkAkMwRqEUSSgAgOkCbCiYKbgm6uh2imtql34+holwVuiv5dt8dtQ8SbdBwcd8x++wfwLQv/+QLI7aCuG7X99n1vOBU6L667zC3N5ODpwhG0b4Qjj3qH7MCwjRBCJEBN7w9KUlCaQjJA7NvHAOH7C3IM3cyv73yQRV7qvG46iLcKo/2ttW/t+xB5nITfgpSyLWCEOIskSbBarVCWJYwxAG6isN61vof4/xGJRCKRyFPlXS7PrtNDa932+UjTFEIIOOeQpimGwyGm0yn6/X50fjwxmlqaBVB477fW2hURLbXWl1mWXSZJshRCrNM03Wmti81mE3rgxpONB0gUQN5ziMifnZ3h9PTUJEliV6uVASBXq5UQQkgikuPxWOZ5rrTWUkqpjDFKSqmEEEoIoZIkUUH4kFJKVQ+VU0SkmFk2QohC4wYhIiHqDs9tRFa4jkYEORA6BFHdO0RK2bpCmmWpcX0EcQSdx90SS7z34nB+NxKrc+Lariv0K+l+ZN3PrxtpFdwn7/q4v+v3ciiAhNGmQoi7+n0Ex8adTo7wuGbjCzTCR6NGh8f5zvIcHB9BCPHeOymlCwKIlNICsERkARhmLpm5klJWzbRk5kprXQKoBoNBVZalTZLE/vGPf3QfffSR/eMf/+iOj4/96ekph3i27/r5PBDoyy+/lIPBQA+Hw7Sqqr73fgBglKbpZDabTX/yk59Mj4+Pp8PhcNzr9XTzv3TfrzvyhAkH+RwamQNN/486/kpUBrKqavFjvwcVBZAXtSDSuEBqJ0gTmQVAMkMRQYmOAIIw6r7Z7nbFjRsN+taRX/dxbQGa35Qdurdv/T91FiN8y1HlO/8NqXVT3LHq7yWCtDugjrnlrtit2zFZuMm14nfLL92hQ54B3wgZnmvXB4MhuP7Imepm5yQlRJaBjK1dO80LdAAg6mXqJukMJm6MK4Rv9z++n3SFjzCCD7j57QQ3iNb6Vo+QyNNCa43RaNRmeSdJAmMMjDFwzr31N9EVLyORSCQSiTws3rUfD+KHcw69Xg/D4RAvXrxoRRBmhpQSSZJgMBhE8eMJIoTwUkqrtS6SJNkmSbJKkmSZJMml1vpKCLEGsCWifDweV9Za99lnn/HZ2dl9v/TIn0EUQB4ATeGZmBmff/65B2BPT0/p1atX9OLFC6qqSlZVJWazmej1eiJNUzkYDKRzThKRSpJEAlBaa6mUksyspJTSey+llFIIIb330hijREMQPYIw0b1eG0luHCDOOeqII9SMzGyXCQJImOmca5dzzpGUEt77VgAJt4UQQbSgO+bditW6S+ToCiNvEz++hzhy+Lg7z5SbmAXuLhNEDADcZE+ycw7deVLKWwKIEMJ3lwnCRxN3xc45FkL4cGmED091g3PXmVoiMgAqa61JkqTKsqwyxpiyLI0QwpycnJiyLC0R+f1+7wH4f/3Xf+WXL1/65nN8bFUBcXZ2JgCIwWCQWGt7+/1+aIwZ53k+tdZOiWiqtZ6ORqPxeDwejEajTEpJoQlOJHJfUBtRRaBg8W6anJMxoLIEihy8z0H7PVAUoH0OLnL4soKwFt7auleIq/uCKAYkAQIEQTgoIN9U9olEU0T/9n4SFOKxmmyn7+PCOFzrtzlAmp1RuzDfoY4cruPbXChvvI5O/NUb9wfh53BV/q5X8ubzh49J4LYIEkQgTwSm2vnhpQKUgqsqSGNbSwlx0/heEFwwgJBqBawgfvjwepsIs4dAt3DdFUHCVErZ9gUxxmC1WrWNK5MkgdY6xhg8AaSUSNO0jbYAgDzP299JiMMKBZK37c67Am4U0iKRSCQSeT/pDgrr7q+7rg/vPay1rUtYKYXBYIDZbIbBYNA+NhxPxuPFpwEzO++9s9aaoii2ZVleM3OIvXotpbzSWl9LKde9Xm+72+3y/X5fXl5e2v/xP/7Ho4mDf4pEAeThEGKx7vpns2dnZ/TXf/3X4uTkRJyfn4vRaCR6vZ7I81z2ej1ZlqWcTqeiqiqplJLGGCmlFNbaIIIIa610znUdIEREZK0VSZJ0XRxUlqVoTjJviSEAyDlHTR5zK5AAgLWWuoSihVIKzTLtsmmatuJIVyQJt4EboaT5DN4adxWWfxvddX5XpJS3voduU63u/UKIVuBohAsglASb20mScIjE6i6bpukt8SM8Rkrpw9Ra295mZi+ldL5Wtlxz2zrnrHPOpmlqjDE2TVMzmUzMZDKxX3/9tZvP58HG5wHwJ5988pg36HR2dibm87mcTqdqt9ulWuteVVXDsizH1tqptXbmnJsy81hK2U+SJEnTNG4rI/dOG68UxI/QA4QZcA5sKqAqgaKoBY88B/Z7UJ4DeQ4qK3hroZwDWwtUFaS1EN61PUDaEwiiWwFQJFod+61RVofFQgriB3dFih9o8/KOLTYdWB1uunTcnvd9n+bOp7zDFhK+p7ftscP9/OYjb1w9AAQBTAJWSEBpeCnhlK77f1gL1wgejV2yyZkkyK4LhByEqF0ijPo7bnIU2z4uD4HuyW13GhwfUkowM/b7PS4vL9uT3slk8kZkVuRxEr5nKSX6/T6898jzHEQEpRS22y3yPEdVVe3voSuCHAofoYASRZBIJBKJRN4vDt0e4fbbxA9rbesGTZIEaZqi1+vdx0uPvAd4770xptput9s8z5fb7fayKIrXAC6VUldSyhUzb5VSe6VU0ev1qjzPba/Xqw36kQdLLOo9Dvjs7AxnZ2f+7//+7/H73/+e/9t/+2++3++LPM89ADcajQQRiSBwVFUllFJCSimKohBKKdGIEiSlFF2hwnvfujaqqqI0TZEkCVVVRUmSgIjIGNNed86RtbYVILTWsNYS1309IIQgay2FyIo8zymM1gyCRmNVpFDcCI9jZiRJEtYXYjHednZKALoCy52ETMg/l+a9tre74kgjZqCqKiilOEkSttbWX1ojgDjnoJTiJreavfe3orOaz5CZmY0xoJt+IUxE7JxjAKyU8lprX5YlG2O81tpba71zzhlj3Gw2s1prt9vtXGiU/uLFC4eO+PHI1Wzx8uVLms/nUkqp5/O5rqqqVxTFsKqqsTFm6pybG2PmVVVNq6oaWWszrvvjRCL3TisihCIdAHgP8h4wFigr+KIAF0UteOQ5OAggZQkUJaS1gLUgY5AUBURZQDkHgZuifdievRkbdVsAuXuZA7oFxb/4E/jz+XOfuytSvHsdByPP/oznItwII2EqtYZQCTjN4HQCpxOwUiBnIdnXoggRJGqRioQACQkSshY3QoG3mbpaBWkdIA9lg0+dCCzgtiASBBDnHDabDcqyxHa7hTEGUkporZGm6X2+/MiPjFIK/X4fz58/R5ZlyLIMzjnked72jOk6RYA3f2Pd65FIJBKJRN4fugMVAuF2qK9472GMaQWQcP1w4Grk6eG9t2VZ5tfX15er1epivV6fO+e+NsacJ0lyKYRYNU3Py6qqzGg0sqPRyH366afR/fHAiQLI46EVQU5PT+n8/JxGoxH3ej1/fn4uPv74Y5JS0n6/F8xM/X6fttutkFJSURSiifehMB0MBiAiyvOc+v0+iqKgPM+p1+shzGv6bwAAGocIiqKgLMtQliUBQLieZRm01qiqisJ9QN28NMsyBGGlO0ozCClpmqKqKmqepxVHDj+Aw8xGY0y7THj8XTRukz/zY693wGVZhtcQXB7QWnMTiQUiQoi0EkKgqqrwWG7eK9I05e56GrEnzGMigtaai6JAcIeUZYk0TZmZuaoqllKylJKFEGyt9czM1lrf6/Xcdrv1k8nESyn98fFxUK+fivhBv/zlL+nVq1dSSqmHw2F6fX3d894PjTHjsixnzDzXWs97vd5iMpnMRqPRWGudElEUQCLvB434Qaj7ftQXAN7XF2vhq6rt+4E8B4qicYQUEFUFbyzYWQhj4YocvqrgrKljtG4913d8ST/8u/zB+SE2bHe5SN7GD/GZ1LY/gtcJvHZwzPDOw1nbCCBJLQII0XGM1CPgWQgIGQQQCa8kPAhEgBSi3ugH8eMBFXjvGu3XjS0IJ7xlWbYDG3q9XnuSnCQJlFLRDfIEEEIgSZJbDo/9fo+qqt5oigrcHbMWnR+RSCQSibxfdGOvALwxOMZ737o8iKgdAGGtxXA4RK/Xg9Y67uOfIMzsnXPeOefzPC+22+12tVotr6+vX2+322+UUhdSytdSyiURbZ1zeb/fr8qytOfn52673fpPP/304Zw4Re4kCiCPCz47O2PuNA7/4osv6Pj42H/44YcAQMvlkqSU9OWXX1KapvSTn/wEVVWR1pqurq7o5OQEy+WydWQcHx/j+vqattstAcBms8FsNsN6vW5vT6dTTKdTrNfrEH3VOjn2+z3G4zHC4wGgK4AAaIsSd8RItevqrBdE1N7u4r3HcDh8Y/5+v6e/xOHxXQivp9/vv7FR3G63t+7v3gbqzxCo3SLd9xnmhVGLw+GQ1+s1ALS3Q2SW956FEDDGwHvP0+mUz8/P2VrLxhheLpf8d3/3dx43cfO3Lo9c/MDZ2Rm9evVKvnjxQhlj0u1220+SZFiW5bSqqrm1dp6m6aLf7x/NZrOjxWIxXywW436/nymlYrUs8l7QbthDHxDnm/grDzgHbwyorMBFCZR1DBbyvHaEFEUtjlgLNP1CtDWoTFX3D/EexL6NU3pMPIRTnG4/kVqZJlghYBgwACwA5xnO1j1A4BzADE9U9/UIBVspIZqpDAIIAE8ASwULBjHdNHV/BKPcQ/RRN+oAAK6urqCUgrUWZVliNpuh3+9HAeQJENzD4ZiKmVEUBbz3UEphv9+jLEsYY9pBKmH6NvEjiiKRSCQSidwfd7mADyOvALRRmIPBoI1Idc5hOBxiOp0iTdO39gGLPF6cc74oCrvf76vdbrfdbDbX19fXl9vt9jzP8/MkSc6zLHudZdmSmTdElJdlWX344Yfmyy+/dP/yL//y6GtmT4EogDxCwj8mM+Ply5e3YsZPT0/xxRdf0MuXL/HrX/+a/v3f/x2///3v6dNPP8VoNAIAms1mrRhxdHSEo6Mj/Pu//3t71ncoNHz00Uf4j//4j1tnhf1+v71urcVyuWzvv7y8/IvOID/44ANcXFzcuY67BJDua7kPdrtde73f7/NqtbpzuSCEdOn3+7xcLgEAWZZx97147zEajWCtvbUh/vjjj/nVq1cAAGMMbzabNlILB4k1T2Ejzsz061//Wvzud7+Ty+VSDwaDlJkHxphJVVUz7/3cGDMfDAbz0Wg0/8lPfrI4Pj6eTafT8WAwSLTWsVoWeS9g5rqHQ3B/oOn/4WsBBMaATQUuyzoOqyzr6KuyBJdl3SS9EUCEcyiZ68baTWQTOW5jmCL3hwfBCIFCSORCoELtEnRVCS8d4CzIO3hmONz0DGEpwUpBSAGSCpAKpBS8IHgpwJLBEHU/F75pR/+QdwLdGKxQ8A4nwpvNBsYY7HY77Ha7Ng4ry7J7ftWRHxOlFHq9Hk5OTpAkCfr9Pr755ps2CiP8dgDcEkGA+vcVnLyRSCQSiUTuh7sanod9dRA/Qo+PNE0xHo/x/PlzDAaDNk49HAMMh8M3kkMijx/nnN/v99Xl5eV2tVqtttvtdZ7nS+/9Uil1pbVeJklynWXZioh2xpjSWmv/z//5P/7rr7/2Z2dn/r7fQ+QvJwogj5iD4nbrDAmiyM9//nMAwG9+8xv61a9+BQD47LPP7lzX7373u7fWxH73u9/h5cuX73wtH330UXv917/+9a113VX4fxf/7//9v7fe97d/+7ffa10/Bv/3//7f9vrV1dX3euynn37KjXvnTr744os35n388cd8enoKAPj888/x2WefvVHfegrCRwMBoIuLC2GMUf1+P2HmHhENjTFTrfVcSnnU7/eP5/P50dHR0fzk5GQym82Go9GoF/rk3PebiESA282fqTsKqnGBeGsbEcQ0U1tft/am6bn3YOdgG9cHULeEsAQknf4ikfsh5BI6EAwRDADjPJxvco49g33j/ggOECHghWgFEKggfkiQFJBSwCsJ5pteLv6OfiMPicMIBODGNRoEkKqqUFUVvPdgZoxGo3aZGIf1dBBCIESsBqdHWZbtbyM4hrojR4GbniBR/IhEIpFI5P44dGAeRl6F+7XW0FpjPB5jOp1isVhgNBq1btAwUEZrHfftTxDvvbfWltvtdrfZbNbr9XoJ4IqIlmmaLrXW10S0ttburLXFfD6v/vmf/9n94z/+o3tCtbNHTxRAnhDv+Mdt55+dnf1IrybyY/GUv9OzszP6/PPPxenpqRyNRqooigRAX0o58t7P0jQ9yrLspN/vn8zn8+PFYjEP4kev14tDQyLvHaH/R9sLJNz2HuR83ePD1sIHG9Neh7Ug6+CdbXuGODBE4yKo8/Hisd37QC2CMBzXsVeefG3f8x4sHNgJwDcChhDwom52zlICWjcuEAmhNaA1ZKrhvIJkD2ZqnERNjxH/MAczHUYRdYvVIe6AmVGWZf1+hcD5+TmA2k0zmUxiHNYTITg8QuY3ESHP81b4CHFYYQTp20SP2BQ9EolEIpEfl7v2u8Gd2RVAtNZI0xSDwQCz2Qyz2QzT6RTD4RD/1VHokQeDc85VxphtWZbXZVleKaWWWuulUupaSrnSWm+SJNlZa0ullGnEj4d5shS5kyiARCKRxwqdnp4SALHZbJTWOrHWZs65oTFm5pw7Ho/Hz4+Pjz94/vz5h9Pp9Hg8Hk+Hw+FAax23jZH3Eu4IH+Ba/GDvo5VGTAAAIABJREFUQY2zA96DrYNvXB/kHNg6sLUQ3rXLgH3t9mgv8djufeEm2sxBUN3kXKBuXC7Yw7MEQHWT89AzhAgsBFipetq4QSjREGkClSb1b0NKcNM3xKOOVHONWPAQ+xscNq8OhesggIT5+/0eX375JXa7HdbrNf7qr/4Kz549Q5qm9/K6I/dDyAU/OTlBlmUYDAb45ptvcHV1hTzPAdyIad2ojbsKMA/1fyYSiUQikYfAXY3Ow/xu74/Q9HyxWOD4+Biz2Qyj0QhZlkWnR6SFiLzWusyybJ1l2bIoikut9ZWUcpkkyTWANRFtpZT5xcWFvbi4cJ988kk8QX5kxCJfJBJ5jNDLly/Fn/70JzUYDJKqqnpFUQwAjJRS0zRN51LKk+l0+mw2mz1bLBZH4/F42u/3R1prJYSIw4Ij7y31QT8gmpMBgboIzkHM8E1zdAbYh2I6g/yN4EGeIdhDNi4QER4beS8gZigwHNfuD0H19+w9wTdfU4ivEkH8kAq+cX+w1kCSAEUKylIIk0IqDZa1o0QQQVDt/CGi2k3yAAu63dfc7QfSjTEKMUer1ap1vMxmMxhj7udFR+6NEIM1Go1aR0iISmNmGGPa0aTBORLEkEC3IBNuP7T/m0gkEolEHgrdyKvudaDu85UkCYbDIWazGRaLBWazGbIsg1IqCiBPHF8f+DvvvTPG7L33ayK6llJeJUlylSTJMkmSlVJq673fb7fb0jlXvXz50sfYq8dJFEAikcij4+zsjABIKaUmosxaO/Dej4ho0uv1Zv1+/yjLsmeLxeLZfD4/Ho/Hs+FwOErTtHffrz0SeRd1MZxA1FzHjStEEOC5cQvUikgrahBqwYQasUMyQzGgmaFR346nCPdPcPdIMBTXnToEAMeNy4MInrjtFcKN+EFCAFVVN7xXCqw1OEkgehlQlpCmB0oc2Lu6KXrzeEEE3xRwH2IvkO4o/XDpNq0mIhhjwMwoiqJtjhmisSJPiyBqhAxw7z2KokBVVQCA3W6HoijgnINzDlLKVjQB3oxe6xZioggSiUQikcgPw12ODwC3mp1LKdHr9TAYDDCfzzGdTjGdTjEYDGLsVQQAwMzOWltVVVUURbEqimLJzJdSykul1FWSJNdSyk2/399tt9ui1+tV//AP/2Dv+3VH/uuIAkgkEnlM0NnZGb148UL2ej19fX3d2263Y+fcxHs/9d7PtdbPF4vFB0dHRx9Op9Pno9Fo3u/3e1LKuD2MPEiIACEITAIkCJB1QZyFAISoY5KImlH/ApIYmggpMzIAKTM0auEklvDuHwGgPm2rv5e6P0s4Aay/SwfAAShJwFkLFhKQFVhreClBjQOEdylElkGUJaAVpBBgAlhKeBJwnUi1hyoHdEWQcLsrgARCc8zY/DwC1GJIr9fDYrGAlBJZluH8/BxFUbQ9Qbq/l7vcIN3fXBTUIpFIJBL5yzgUPsKUmeGca129UkporTGZTHB0dISjoyNMJhOkaRqP8SItzjmT5/luvV4vd7vdN9vt9quyLL+21p4rpV4DWKVpupVSFtZas1wuY+TVIycW/CKRyGOAGteHOD09FcvlUq3X64yIht77KYAZMy+stUda62e9Xu/5fD5/Ph6PjweDwURKqWPsVeShIohAaApzjehBzZSbeUwESQSJesefAsjAyJiRAJCIAsj7QvgeBOrG9OFUsDkNBDPBeYYBQI5giOCErB0gUoFJwDcN0CnLgKKAKEtQogF10wNEoomLIgKY4W89z8PirgK0EOLWyXMoZgdXSFEUyPO8HeUfT5ifFkIIpGmKyWSCJEmglIK1Ftvtti2yaK1vOUBCEeZQYIviRyQSiUQifz53xUuGqfe+vYQBL1prDIdDLBYLPHv2DIvFot2XR0fmk4aZmX1Dnuf5drtdXV1dXazX6z/t9/uviOhP3vsLKeWVEGJtrd2Nx+NiNpsZpVQUQB45UQCJRCIPHTo7O6OvvvpK/s3f/I0oikI555I0TXtFUQy99xNr7dw5t/DeH3nvj5RS816vN+33+6M0Tfv3/QYike8KgW7FWlEzT9BNU2yEBr5BEGkaZksiKAISAAkzUgBJ4zKgWMB7P+g4Mt4eScZwEJDe1c4eJ2CsqaOtqqpudF6W8FrXwkdZgYoSIk0AreGFhBPBDdT0AUETq9Y8PzPXv6UHyGED63AiHBpleu+x3++x2WygtUav10OWZVEAeWIQEZRSbRwWM2O/32O1WkFKCedcO997j6qq4Jy7tY7Dkaqx6BKJRCKRyPenO5DlsMl5iL0C6sELSZJgNBq1kVfT6RSj0Sj2+4gEp5C31pqyLM1ut9us1+vr6+vr1+v1+iLP84skSV5nWXaltV4B2AohCgBVr9ezv/rVr6IA8siJAkgkEnno0FdffSX/7u/+TnrvNTMng8Eg2263I+fcxBgzc87NrbULY8yiqqppVVUD55xm5nikFHl4NCP2D4tt1BE/fCgCAwDqorYC17FX7JGwh2aPWPJ9mBAYkoHUOwjUDc2NEDCigpcSXGpQYsBFAZQlqKpqIUTrOgoNBEkCUgj49ndUB2FxGH13b+/uL+ewGB1isZgZZVni4uIC1lrsdjscHx9jPp+3TbEjTw8hBLIsw9HREYQQyPMczAwpJYqiwHa7xdXVFfI8h7W2fUy32BLEtfgbikQikUjk+9Pdfwbxoxt7pZRCmqaYz+c4Pj7GbDbDfD5HmqZx3xsJsLXWbrfbfLVabVar1eVut7vY7/eXTe+PpVJqZa3dMPOWiIo0Tcvz83MLwH/22Wd8dnZ23+8h8l9IFEAikchDhn7+85+LDz74QHrvtbU2TdM0K8tywMxj59zUObdg5iMiOkqS5EhKOQUwBNq2B5HIg6MbjQRBbXZVE4YF0dxmqu8TqHf4CTPSRgBRTePzeMrw8AiN0sl7CFiQA9gIeCHBxgDG1JFYTWN0FCWQJBBJAiEllFRgr+A9wxPXMWmN68OFUe0P0AVylygYIouklPDeoyxLWGtRVRXKsmxPqENE1mFhO/L46cZhZVkGa237u9lsNri8vERZlnDO3YrAuktoi0QikUgk8udz6P4IgwuSJMFgMMDx8TGeP3+O2WyGNE2RJEnc/0YA1L8dY4zN83x/eXl5vVqtXu/3+9fe+9dEdJWm6VIIsdJab7TWe+dcAcCMRiP3q1/9yv/DP/zDQx7/FfkORAEkEok8WF6+fCk++eQTcXp6qpbLZQqg770fWGvHzDx3zh1574+11idpmh6naXo8nU7ng8FgpJQKrQ8ikQfETUYuEdoCNXX7gAQ9pBVFao1EgqHA0FxfYon34XITk8Ug9oCz8CAw1U3vvVKA1kBZgfMc1MvqHiCJrgv8UkE0fS+UJIBvmq23MQQP7GSye/J7V4E6OECcc6iqCtZaOOeQZVl7X7/fR5Zl8WT6iRHyxJVS6Pdvp2ImSQIAKMsSRITtdgtjTFucORRADvuBxGisSCQSiURu0903hut39f0AACklkiTBeDzGYrHA0dERFosFxuPxrajTSAT1qYwxxux3u91ytVpdFEXxTZIk36RpepEkyRWAVZIkW+dcvt1uq9FoZD799FP3s5/9LMZfPQGiABKJRB4q9N//+38XANR6vU6EEJlzbrjf7yfe+6lz7tg5d8zMJ2maHi8Wi+OTk5Oj4+Pj6Xw+H2ZZliilYg048uDgw2lozHtjBGnjr0IIFiH0lrjpMQGOg1weLJ3vLrhBEu8AZyAtwRgNZypwWYKLElwUIJ0AOgFJCdE4HaRS8FKAhYBD3QidOr+jh/oLOSxChwis7v0hDuv169ew1qIsyzZSQUoJpeIh8lPjrkJKmqYYj8etWLZcLrFarZDneVuc6fadAe4u5sQCTSQSiUQit/eRYdo9bgvihzEGSilkWdYeny0WC0ynU6RpGt26kbtgInJSykIIsZZSXkkpL7IsO9dav07TdOm93wIoqqoyeZ7bP/zhDz6KH0+HeHYXiUQeIuKXv/wl7XY7WVWVJqLMe9+31o6EEFPv/RGAYynliZTyeDAYHC8Wi6O/+qu/ms/n8+FwOMySJFFSynjk9D04bPgauU9CnwauG6CjLlYLOlgiCCPMtVvgR3+dkf9qCIBkD/IMcoCwBG8r+CYCi8sCfp8DSoMSDdISpBSkUmBr4aWAByCJwKL+HXX/ux/Df3qILQp9HcLoQmstrq+vURRFO8I/SZJW/JBSxsL1E0cpheFwCK010jSFlBLGmDYOKxAKOG/7vUQRJBKJRCJPne7AgDDtiiDdC1C7MIfDIU5OTnB0dNTGXsVBKpEODIAbLBEVSqltkiTXWusrY8ylUupSKXXV7/dXZVnul8tlWZalAeB+8YtfRPHjCRG3HJFI5EFxdnYmXrx4IVFvv1IAvTzPh9baifd+JoRYADgSQhwPh8PjLMuOFovFfLFYTKbT6Wg8HvfSNNVCCFCsRkQeMoeV6g6tywOA9AzJHtp7SM8QUbx6VITvmpgB78HOQjoHaw1cVcKXJVyRg7WqY7CUAksJSAVqCvwiAYSgpqF67RvyQG0HYX7QIkh3dH7oAyJlnX4YeoGESKNer4c0TcHMGI1GyLKs7QsSeZoopSClhNYaAOCcQ57nICJsNptWDAlxWO+KxQrTeOgRiUQikafE4SCAw/1icFR679tBK4PBAMPhENPpFLPZDLPZDKPRKPZqixzC3nvnnKuMMbuyLK+rqloCuJJSXqVpukyS5DrLsnWWZbvJZFI458zFxUUQPx7yaU7kexIFkEgk8hCgs7OzcNSkUMdeZczcBzD03k+ttTPv/bFz7lhrfTIYDJ4tFotnR0dHJ7PZbDqbzUaj0Sg6PyKPh6awS6A7D90E6qJ44iy0tdDGQHsH4ugEeVSEoioapw8zYG3t7qgquKIApISQEug4GuqeIQC8h2CG0ApCSQgCmKhuiO651kDu79394IQ4rCCEhF4geZ7j4uICzjnsdjucnJxgsVig3+/HE+0nTBDQhBDIsgyTyQTM3PaKubq6Qp7nsNbeWvZd64tCSCQSiUSeAu9KDwhuXADtsZi1tm12PpvNMJ/PMZ/PMZ1O0ev12sEIkUiAmdk5V5Zludrv9xf7/f7r7Xb7n9bacwBXQoiV936rtd4bY8rdbmdHo5H7+c9/HsWPJ0gUQCKRyHsNMxMA+vzzzwUA8eLFC+WcS4UQfefcuKqqsTFm7pxbeO+PmfmEmZ+laXoynU6PP/jgg/l0Oh31+/0sTVMlhIgVh8gjoDleI2pjsEIxjToX6T20c8icg3YOoil2Rx4rtQsE3oGcBWwFVxaAFPBS1AKIqBulQwgwUS2GNVMBQChZ/7qI4IP48QCbogfeFj0UXCBa6/ake7lcYr/fI8/ztiF2lmU/9kuOvKdordHv99seMVJKFEWBqqpa50eIWjt0gQTuavwaiUQikchj5S73RxA/QpxkOA6z1iJNUwwGA5ycnODk5CSKH5G74EZQY++9Ncbk+/1+eXl5+dVut/tyt9v9Z1VVF0S0BLCRUu6rqipXq5X98MMP3b/927/5n/3sZ/GE+AkSBZBIJPK+QmdnZ/T555+L09NTcXp6KjebjVJKJVVV9fI8HzPzFMDUOXfEzEda65Msy056vd7J0dHR0WKxmE4mk+FoNOqlaaqISMSRvJHHQ2dUVZOHdau5ufcQAKR3EM5BeR/dH4+c0Oheeg/VOEC8kHBCAEK0DhBqBBASBCgBEgJCEFgQpBB1LxBmSEFwTWH3oZ4ldEfbH14XQrRCiHMOZVnCGAOtNfI8b6ONIhEAEELcyh733mO9XrcxWOFirYWUsnWC3NXk9bAJbCQSiUQij4Xuvu2uhudB/AjHWSGmNEkSTCYTzOfztuH5aDS6tU+NRHATe2WMMfs8z5f7/f58u91+tVqtvq6q6hshxCWAtVJqlyRJXpZl5Zyz5+fn/tWrVw/1tCbyFxIFkEgk8l5ydnZGL168kEmSSADKGKO998l+v+855wbMPGlcH3NjzJGU8ijLspMm8up4Pp/PZrPZeDAYhNgred/vKRL5obhp/9E5fuNOUxAOggiDGHXEEfONOBJ5nDTfs/YWbOqIK0MClgieCNyIHkRUix5SALIWR6Sue4OwFJAk694f3EQA4eF6xN/Wg6EbgxXu656UhxPyWJyOBA7jsEajEY6OjiCEgFIKm80G+/0e1loAuNV3ptuLJhB/X5FIJBJ57HSPwcKxVYi86sZe9Xo9TCYTLBYLHB8fYzqdot/vI0mSe34HkfcN7z1ba01RFJvdbnddFMU3m83m6/1+/7Vz7k/OuddCiKW1dqOU2u/3+9IYY3772986AP7s7OyhntZE/kKiABKJRN5HCIDY7XaqLEtdVVWilEq89z1mHjDzyDk3d84dWWuPggDS6/WOT05OTl68eHE0mUzGg8Egy7JMSSljhSHyKHnj6I1vnCD09qUijxQCIJmROAfB9W0PgiWCI7oVgRXED1ISUAqUJLUYoGQdrUYEyXUM1kPfgB4WnsO8w7iiEK+gtYbs9EuJRA5RSmEwGODZs2fIsgxZlrW9ZIwxt5b9tlgsIIohkUgkEnk8dN0e3UbnQQQJg02MMTDGIE1TjEYjfPDBBzg+PsZ8PsdgMIixV5E7YWZfVVW52Wyur66uvtlut/+Z5/lXzrk/AbjQWl8qpVZa641zbr9araqf/vSn5uzszIVV3Ofrj9wfUQCJRCLvE/Ty5Usxm83EeDxWRJT2er3UWtvz3veIaOi9H1trJ1VVLYQQx0qpxXA4PBoOh0cnJyfHi8ViPpvNxuPxuK+U0lJKolhViDxqOs6PyJMmNEIPUWfOAcIKcNU4QA4isCAESClIpSHSFEIpkFKgpj8IA3U0VugVgof7S7ur70KIwfLet6P4gfokPc9zbDYbKKXa0YlKqRjBEAGAViDrCmV5nsN7D6112yOkm21+GKd2VwxWFEIikUgk8tDoOmzvIuz/iAhpmrbHUmH/GByVJycnWCwWGA6HkFIiBjhEAszsvffeWmurqsr3+/1yvV5frFarr1er1dfOua+11t9orV8rpa6ZeVsUxT5JknI4HJo//OEPsel5JAogkUjkvYF++ctfilevXsnxeCwHg0EihEgB9LXWA2YeGmOmzrmpMWbmvV8Q0XG/31/M5/Oj+Xw+Pz4+ns/n89FwOMzSNNVCiHjUFHkSvBlSxG9GZEUeP+EEFKgb3hM1zdAFICpwKWsxo+kHwlJBJgmQphBlD1CqvjSiBxPBoRZCuqXbh/qruisKq+sECSfk3nvsdju8fv26bco5mUwghIgCSAQAWvFDSol+vw/vPYqigJQS+/2+FUaqqsJut8Nut2sLQEHk6Oajd6dRBIlEIpHIQ+Ft4kc3WjS4P0LU1Wg0gta6HSTQ7/fbnh/9fh9pmt7HW4m8xzCzt9aaPM/3u91us91uL7fb7ev9fn9hjDn33l+kaXrpvb/23m+klPtnz57lVVVV//t//2/32WefxaZ+kSiARCKR+4eZ6fPPP6dXr17J09NT+ac//UlrrZOyLHsABlLKsbV2wsxHzrk5gLlzbqG1Ps6ybHFycrL44IMPprPZbNLv91OttY6uj8iTgPmgGl27QaL4EQEAeAa8B6wDkwGLOt6KpICXAkJKIG0EkH4PlGgIYwCl4IWDFAKSASZAoBZBCM3J7gPcxHYLzOF2mBccICGW4fr6GkVRtD0dtNbtyP5IpIvWGoPBACcnJxiPxzDGQEoJay222y0uLi5gjGldIEKIN2LZYkP0SCQSiTw0DuNFD+cHAcRaCyEEpJSYTCZ48eIFBoNBe9yltUav18NwOIzHWZE7cc75qqqq6+vrzfX19evVavVNED6UUpdEdOW9vxZCrJIk2SVJUlZVZZIksQA8EcUT40gUQCKRyL1AzIzPP/+cAIgvvvhCjMdjqZTS5+fnOk3TZLvd9qWUI2PMGMAUwNRaeyyEmGutF1rrxXg8Xszn89lisZhOp9PxZDLpKaWUlFJEASQSiTx1BBjSeyg4OCI4aeAFgcs6+opVAZQZqCxBeQGRJPBKQ0gJSQQWElIIeAZEs0n16AgJ9/je/lzuKjIHIaTbHL0oClRVBaDu95BlGYiobcgppYxukAiAWjxLkgREhCzL2t9YiE4LGecAUJYlnHNviB9h2hXn3lZYikQikUjkvugeR911un3Y6yPEXmmtMZlMMJ1OMZ/Pb7lAgjgS4iMjEaBudt44P3xRFMVut9ut1+vr6+vry81mcwHgQkp5KaVcCiHWRLQlor0Qonj27Jn56KOPLAD/s5/9LB5QRQAAcesSiUR+TAgAnZ2d0W9+8xt5enoqlVJ6Op3qwWCQaq17AAbe+1ETcxUanR9XVXXsnDshopM0TY/n8/nxycnJ0bNnz2ZHR0fj6XTa7/f7qWyafuDh9+29d4qiwG63w3q9RlEUbzR2DUSt6ceBDi/MEMwQxkBUFWi/gyhKoChAlYEoS8iqgi5LKGOgnHv3E0QeF00Pj3DETwBAoo22oiYKS0gJqVTT30JCKHXTH0TWkVkgAgR11vRm6NpD4a6R9nf1YQjRV+EEPjhDALQn6vEkPQKgFc6UUkiSBGmatj1jukWicN1ae0sEOYzDuut6dIdEIpFI5L55V6+Pw8ircFFKYTAYtMJHaHI+Go3Q6/XafabW+lZfrUjEe++NMXa325Wr1Wq3Wq1W19fX5+v1+pvNZvMnIvpGKXWhtb7s9XpXSZKsyrLMy7Ksdrud++ijj1x0fkS6RAdIJBL5MSAAODs7o9PTU1oulyJJEglADYdDvdvtEiJKrLUDAANjzMg5N3bOTZl5aq2dNZeFlHKWpuns+fPn0xcvXkzn8/mg3+8nWmsVD5h+POLo1PcDCn/aK3dNI08RQj3KJWUPwYDyAJwFWwGrFNgYoKpAVQUUBXi/B7QG6cYBIgVYSkhRN08H40ZUYQY3P6+HWJg9FDzCCMVub4bQwNpai9VqhbIosd/tURQFlFLQWiNJknt+J5H3GSEEsizDdDptxREhBIqiQFmW8N63v7PAXS6Qh/b/FYlEIpHHR3dfdbhvCq6P0NMjXMLx1HQ6xbNnz1rhI8uy6KKNfCvOOZ/nub26usqvrq7W19fXS2PMVVVVl1LKSyK6ArDUWq+EEDspZemcs1999ZX/x3/8xxh7FXmDKIBEIpH/Kujs7CwcGYkXL15QWZbiyy+/FGmaSuecLopCp2maElEGINvv96PG/TERQkyTJJlrrecApsw8McZM+/3+ZDabjReLxXixWAzG43FPKSWklPEoKvKkuFUSYz6QO6IIEqn7dmgAghlgD+MdrPdw1oKUAowBl7VrCGkKJAkoSUBSNiKIAisFOHcjfjQOEg8GNb1AHmKR9m1OEADtCMQwSr8sS+T7HAyGlBKDwQAA2oaeMQ4rcheh8NPv91u3kDEG+/0ezIyqqm4Vje5yJR06k6IoEolEIpEfk+/S56Mrfnhf95qWUiLLMozHY8xmM8znc8xmM2RZBq11PG6K3In3nr333lrr8zwvt9ttvl6v18vlcrlery8BXHrvL4UQl0S0FEKsAGyZOffem5/+9Kf2f/2v/+XwMI3qkf9iogASiUR+aAgAvfz/7J3Jjhxndv3PN0ZEZuRUA0V2C+i/G4YXbHilhgHDMMBe2vDKgPwWfgaVXsIvoW2vvGJvG9CyBcNoCDYgi2TNmZEZ0zfc/yIyglmpIlukKA7F+wMSOVZWJRkZEd89957z+ed9X7r81a9+Jdu2lePxWDVNozebjUmSxAJIQgipEGIkhBg552bbyY9FmqaL0Wh0NJ1Oj4wxMynltG3bPE3T8XQ6Hc/n83Ge59loNOIWXOajZr8MtmuTxXzEbEWx/hKIoGOEDB4yKMS2hZASom07EaSqQEqBjOkEEK0BrUFGgaQApEQUAlHKwQ2rt9j6UIuxLxNBelsj7z2882jbFsWqGPJA+sU+dzIyL0IIAb21l+snPZqmQV3XEEJgvV6jrmt47wcP9NveY7/4JKXkCUyGYRjmrbB/HNq/vWt95b0H0B2nRqMR8jzH4eEhFosFZrMZh5wzf5EYY2zbNpRl2RZFURVFUVxfX18XRXG52WzOpZQX1toLpdQlgGsAqzRN1yGE+vvvv/f/8A//EAAQT38wt8F7H4Zh3iR9xod8+PChBKDOzs5U27YqTVN9eXlphRDGWpt471MpZdo0zVhrPY4x5jHGufd+7r1fjMfjg8Vice/TTz+9l+f5LE3TsXMuUUoZa63J89xaa7nixHyUvLzc3C9UeAqEeY6gbmJDxgjhfVdEbVtAawitEaUEhIDQGkKp51MgursNKSG34ocUEkA3CUJ43gGID1AIuU38ADAUo5VSiDrCwMAHj9VyBe88iqJAuanwy1/+AlJKGGPe+t/OfDj0QekHBweDH/r5+TnOzs7Qti1CCN33S8rBhm03A6R/D+DlNiQMwzAM81N50bGlFzsADBkfu7kf3nsopZAkCY6OjnDv3j0cHR1hOp0iyzJuFmH+It77WJZl++TJk8319fVytVpdN01zTkRPrbWnQohTpdT51v7qGsAqhFAqperj42MHgK2vmBfCAgjDMD+VId/j8ePH8m/+5m/Er371KwVAbzYbvVgsdAjBrNfrJEmSBEDStm0WQshCCGNjTJ5l2SRJkhmAuXNu5pybLRaLg8VicbRYLI6n0+kky7IsxqjkFmOM1FrzWRTD9NxaA+PCGNMh0FlhqRhhQkB0DgAg2xZCKUQhumtjIY3pLLK0hjQGUBJKCCitEYSAEgIkuih0KQRib83zbj/iT2J3sS+lBMXYhcFjx+Yhdh38bduCiJCkKQ6PDodwdIZ5EUIIGGMGW6x+umjXDqvvit0tKvXb1m32WD0sgjAMwzBvgr8kfOxegO58qbd47HPTrLXI8xwHBwc4OjrC0dERrLXQWvOxivmLbCdA3Hq9Xl9fXy+Xy+WFEOJMSnlqjDkVQpwrpS6ttUujnQl2AAAgAElEQVTv/bqu6yqE0Dx48MD/53/+Z/zd7373IS9HmJ8ZFkAYhnlVhjOXPuOjDzb/13/9V3l5ealijKqqKtu2rQ0hWKWUJaIsxpiFEEYhhLH3fiylzI0x0/F4PJ/NZnOt9YKIJk3TTPI8n83n88VkMllMp9NRmqbpu/vIDPM+82LTK7bDYnrE1gLLQEAgoHNopudFfgBRKcBYCGNAW/FDWAvS22kQIbpwdJKQAISU8Nv3J9AHOwVyK0JAbq+VUpBCwjmHtm27YrUxqKoKzjmEEN/1X8u85+zaYfXTQs45VFUFrfXQNeu9h3MOdV3DOffSDJD++jabLIZhGIZ5VXYFit1jze5jvTivlBpyrnqrx10B5PDwEPP5HJPJhIUP5kdDRDHG6Oq63mw2m+uiKC6SJDnNsuxZkiSnSqnzGOO1EKIgonI8HtfW2vb3v/99PDk54RNy5qWwAMIwzI/hB6LHn/70JwFAPHjwQAAQm81GJUmifvWrX2mllPXeJ9baNISQOOcyIcQ4xjiJMeYhhAkR5THGqdZ6MZ/PDz/99NOj0Wg0k1KOnXOJtTbNsmyU53mitVbv6oMzt8PFFob5cBDYBqITQcSACAJRBMWAAEIAwQkBUgpBm07w0ArCmG4KREmQklDbTj+SBJISgQApbmaBfKh7ht3sj939mxASSgpEEaFJD0KP0RpGa0gpICUv7Jkfj5QSSZJgNpsBAJqmGSyw6rrGarXCxcUFQgiDn/q+HdbLQmm50MQwDMO8CvtiO3DzfGg35yPGOAggSZLg+Ph4yEMjIiilYK3FfD4H9y8yr4qUMmqt2zRN11mWXVdVdZam6VNjzFNr7SkRraSUq7quq+l02jjn/H/8x3/QV1999aEuQZi3CAsgDMPsMoQGnJyc4E9/+pP4zW9+I77//nvx2Wef4cmTJ+Lg4EBMJhMxnU5FCEFqreX//d//KWutAmCIyJRlmSqlshhjFmPMiGjsnJvEGKfOuakQYpokySRJkvlisVjM5/Ojg4OD4zzPJ8aYJMaohBBKb5FsGMowDPOTkAA0CIoIFAlABEUBB0ILwAuBqBSi1iDT2V9BayitQUpCbjNBtNKgbSYIUQRBDgLIXVh53BQ/elEEENhaPIAAwhBq7bfd+mmSdFMyW3sjhnkRvR1WnudIkuRGCPp6vYbWGm3b3rDCui0I/UXvDbAQwjAMw/xldicJ+/u7z+0KH7vHIq01sizDdDrF8fExFosF8jwf3q+fduytHxnmZRBRJKIQYwwhhA2AlTHmKk3T8zRNT40xz6y1z4wx51LKcr1eV0mS1HVduzzPw1dffRVxN5YhzM8MCyAM85FDRAIAvvzyS/Hw4UMBAN98840AIP/xH/9RTCYT8eDBA5llmXj48KF4+vSpBCCttWo0GknnnM7zXAEwzjlb13USY8ycc2MhxCiEMOqnPrz3MwAzY8x0NBpNp9NpL4Ac5Hl+mOf52HCSLMMwzJuFCAKA2rk/IIDgBdAqBKVAxkDUNeJ2+kNYC6E1SBsIbSC0g9YahIBuOI9AAoh4rqDfCSssomEltVsc2M0J8d5jvV4jTVMoKZGNRrDWsgDC/EV665D97lhjDEIIqKpqKDjVdY0QAkIIEEJ0GTV7HbpcYGIYhmFeh93jye79fQGkPwZprZEkCabTKRaLBebzOQ4ODpDn+Tv7DMyHDRGFEELjnKucc1cxxnOl1LnW+jxJknOt9UWSJJdpmi6bpmmm02mzXq/bqqr8119/zeIH86NhAYRhPlJ64QOA+Oqrr8SDBw8kAJHnuXj48KE8OztTs9lMOufkYrGQANRms1Gz2UxtRQ+tlNJCCFtVlSWiBEDivc+IKAshjEMI4xjjmIjG3vtJCGGitZ6Mx+PJ4eHh9Be/+MX86OhoMpvN8jRNrVKKV/AM8wrwF4b5yRCASEAIgA+Ac6C2RaxrCG0QywpSG0AbSGugjUHQ+rnllRKDADJMgdyFYqwQnVDU23rthaSHGLDZbPDs2TO0bYuyLHHvk08gpQTr+MzrorXGZDJBjBFJkiBJEpyfn6MoCnjvB3FtX2S7TQTp78cYWSBhGIZhANw8Xrzo2LArfHjvh+skSTAajXB0dISDgwMcHh5iMpnweQ/zk4gxuqZpis1mc7bZbJ6t1+snm83muxDCU2vtuVLq2hizJqJKKeXatnVKqfD5558HAHRycvKuPwLzgcACCMN8ZGyFj+Hy1VdfyTzPxaeffiq/++47dXl5KVerldJaq6qqlJRShRBUVVXGe6+11loIYYjINk1jnXMJgCSEkMUYR1rrkRBinKZpL3yMQwgj733uvR9prcej0ShfLBaTe/fuzQ4ODkaj0cgaY4wQgttm32M49+M9g2ho5CeibVf/oGu+q7+K+cAQRBAxQoQA6T1C24KaBlAaURsIYxG1htQaMrGAsYBWg9ARBRAhIYVAxE4oM+7APmMrgog+KH5bNJBSgmLchqC3cM4NhQGlFLTWkFJCSsmFZ+aV6G1FdrejsizRNA2ccwAwTIb02yLwwyLWrnc7b4MMwzDMvt3V7mMAbrVclFJCa40QAogI1lpMJhPcu3dvCDlPkgRac1mReWUidUTnXFXX9fVqtXqyXC7/b71ef9+27ZMQwqm19lIptXLOlUmS1MvlMiilQpZl4csvv6STk5MPfLHBvE14T8UwHwlEJL788kvx+PFjeXZ2Jo+Pj+V6vZZJkqimadR3330n67rWVVUpItJt22pjjG7bVnvvNQATQrDee+O9TwAkABIiSmOMaQhhrLUeG2PyyWQyTZJkorUeO+eyEELqvc9CCImUMp3P56Ojo6PxwcFBPplMEmOM4gU6w7wKvYbZ39u9z98l5scjQJAUYYIHOQcohagUSCmQ1t1FyS4M3VoIY7qsi63mpkSCAHSPbRfWAdutcC9Q/ENiKArsWAz1FyllZwfhPZqmHgoDaZoOhecsy2Ct5a5I5pXobbHSNIVSnWndZrMZvkdt2w7h6L0V1u52CfzQFutD/Q4yDMMwP53d40QvcOyuu2OMP7jdZ1X1No1EBO89xuMxDg4OcHBwgMVigclkwiI781qEEGIIwTnnmrqur9fr9en19fX319fX3xVF8b219tRae+G9vwJQKKXKxWLRpGlK3377bfzjH/9IJycn8S/+IobZgQUQhvkIICL5+PFj+Xd/93dqK34o770qisJorXXbtto5p0MI2ntvYozae29CCMZ7b4QQRghhpJQ2hJDEGBPvfSqESGKMGYA0xjgej8eTNE2nn3zyyWI+n8+zLBuHEEyM0WyFEyOlNGmamvl8nqRpapRSUvCZE8O8PlzbYn4Cggg6RiQAZPBonYPTBtE5xKYBlILUussE2QogtB3WEwCElJBGQ0Igqk6Kk0IgbnNHgA9zE31REXmwwRISQonBIqIsSzx79gx1XWNTljg+PsZ8PmcBhHll+m3MGIPxeIx79+4NhajLy0usVqtBANm93JhQ2hM9xAcsRjIMwzCvR7/f3xU2du/v5330j1trkec5Dg8Pkabp0PiRJAkmkwkmkwmstSx+MK9NjNHVdb3ZbDarzWZzulqtnlVV9cx7fyalPCeiSyJajkajAkC1Xq/dn/70p/D555/TZ599RkIIPqlhXhkWQBjmjnNyciK//vprBUCt12u9WCzUer02bduaJElsXdfWe28BmBijiTHatm0tEVkppdVa2yRJDBElQggbY0xCCInWOiWiNISQElFGRKM0TSej0Wg2m82Ojo+P55PJZExEkohkjFESkQQgpZQqSRJlrVUsfjDM69OFTQMQzxcv/IViXgUJQBNBxggZPCgoRO8QW4coOwGEtIZUCtAGQuvO+grb7U129ldKSpCUAASIYieIPE9F/yBzQW47PA2PSQCx69jvg6qbtkVZVaibBlrrYQKE7bCY10FrjfF4DCklrLWw1qJtW1RVhaZpBrFD7li07Xf37gp4+7YnDMMwzN1kt2njRROBveCxK3wQEaSUg9BxfHyM2WwGYwyICFprGGOQJAk3eDCvCm23v0hE1LZtXdf16urq6my9Xj8tiuKJc+40xngupbwUQlwLIVaTyWRdFEVdVZX/t3/7t37ig09imNeCBRCGucMQkXj8+LE8PDxUdV2b6XRq2ra1UsokTdOkaZpMSpkSUeacS5xzlogSIkpCCKnWOplMJul0Ok3TNLVSShtjtN57G0JIdi5pjDHL83y8WCwms9nsYDqdTvM8z3bD1vu/abtoF1ve4b8Qw3zAiOfFrd1vEYsgzKsgACgAkggUI3QIaL0HtS1ICAQhIYREEAJSbIutBNB20YxtYV9KASUNoLosmgBAEhDxvLvwQxRB9rlRSJaAhEQIoQsIbdrh+TzPkSQJpJRI0xTGGC4WMK+ElBLGGCilhiLWZrOB937IBwG6Tl7nHJxzCCFACDH8zL7f+64wwiIIwzDM3eK27Kfd/f2u6NHf7m08+2NOlmWYzWZYLBY4ODjAZDJBkiTDa3rxndfwzKuw3eZ8jNE559qmaa7Ksjxbr9ffF0Xx/Xq9fiKEOAVwYYy5jjEWADZZltWnp6fu888/92Dhg/mJsADCMHeYr776Sv7mN7+RTdOYNE0T51wKIF2v1+MQwjiEkAMYK6Vy730WY8ycc2kvaFhrRwcHB6Nf/vKXeZ7nqdbaxBh1jFH11lYxRt3fttYmWZZl8/l8nCRJppSy7/rfgPnp8Anu+whtcz/QFaOpa0jvpRAubDE/mn6xjOeB6PAekA5x+zQRASFARAJiBNoW0jsghiEnQ2kNoVS3XXYbI4LottJeFLhLW+VuV6WQEhKAkAIhBFRVhdPTs+H2wcEB5vM5tNa8P2V+NLvZHmmaYjqdwjmHJElQ1zWk7MS3uq5xeXmJ5XIJ7/2wbSqlXlik2u8O3p8QYRiGYT4s9qc79okx3rj0eVK9IJKm6WC7eHh4iMPDQ+R5PjRxMMxPhEIIrmmaYr1eL8uyfFoUxdOmab4LITwB8L1S6lRrfRljXBlj1iGE+n//93/dP/3TP7H4wbwRWABhmDvM8fGxWC6XCoABkEgps6ZpxsaYSYxxKqWcCSFmIYQZgJEQYiyEGEkpMynlOE3TcZ7nk4ODg+lsNsuSJNFbSyuxtbVSAESMUQKQQgitlNJJkhittXqnH555o+yG5zHvlh+UqIb88+dR6P3/Ev9/Ma+CADqBwwcI4QAihLjtEgwBFGMnhHgPSRGdp6GCMgYySTqbLCFAkCAhQCDQzfGkD3oKZBByqJtyEUIiUuwyF4DBIsI5h6urK7Rti6ZpBzsJa+2NznyG+bForZFlGY6OjjCdTgeho21bLJdLOOeGsPQQwo2ffdnUx774wUIIwzDMh8eLzvf3Jz/6aY/dKZB+clBrjel0ivv37+Pw8HCY/OinDRnmNehtryjGGJxzdVmWq6urq2fr9fq7qqq+d859p5R6muf5qVLqKsZYENE6z/O6qqr27OzMA4ic+cG8CVgAYZg7zGQyERcXFzLLMhVCMMYYK4RIiWgkpcyllDOl1FxrvQgh5EqpPE3TsRBinCTJ5PDwcDybzSbj8XiS53lijNG3WVrt3O9traSUklfQDPOm6YtUMYJ2rIW2+sfzl4HFD+Y1IIKkCB0DYpAIAAIBEdvOQdpudUTQSgJKQ1oLkaYQ1gJSQgkgKgWlOlEAQm4zQ9CJIx+wCHLTUmI7eSVFN0SztQiLkRBjgHP1UEzOsgzGdGGhaZrCWsvTIMwr0eeAaK1vCBxt2wlsm80GVVUNeTR9oasvcvUFrN1mhpdm3DAMwzAfBLcJ2f39PttjV/wQQiBJEmitbwggk8kEi8UCi8UCs9kMSZIMk4QM8zpsxbYQY3Rt29ZlWS6LorgoiuLZdvrjSZIkT40xZ1LKyzRNCyIqpZR1URQtgD73gxe1zBuBBRCGubsIALDWCmutVErJEILSWusYo1VKJTHGTAgxVkqNlVI5gInWejIejyfT6XQ6n8/zw8PDUZZlmVLKKqV4quMjpT+ZZt4PhBAQEMM1EQAiEJ7nf3AZi3lVBAiKCDYGkN8umIkQ+m5BAHFreRWNgTQWcZMAWwFEKg0CoK0FQNtQdAK2evgggryzT/hm6UWQ/k73nYwQQoIoDF35FxcXICJ477BYLDCdTiGlBB9SmR/Lrh2W1s+Xb0opeO9xdHSEGCOMMVgul8NUCIDBDqsvZEkpbxTIWPRgGIb5sNgXsfdzPnanAXvLK+89lFLDpEee57DWIsYIIQRGo9Fge8Uh58ybgIgoxuiqqiqLoliWZXm+Xq+flWX5rG3bU+fceZIkF0KI69lsViilysvLyybLMjeZTMLvf/97Fj+YNwoLIAxzh/n2229FkiRiPB4L55wEoJRSSnerZxNjNERkQwipUiqVUmZ5no+Ojo7ye/fuzWaz2Wg0Gtksy4xSilfIHyksfLxn9BMfQ9g5DQ31wyQIf1uZ10ACMBQhibpMCyJ4AAEYrkkICKVAdY1oLXSaQVQ1hE0glIIWAkFKkFDDAt2TQOzFuQ98CqTntuIDgKFTshc3mqbBxcU5qqpEXXcd+kmSIEmSt/9HM3cOKeVgjZWmKUaj0TARUtf1MAWitUaMcRBBbhPf2P6KYRjm/WdXvN615uwnPnqLq91JwD7vw1qL0WiExWKB+/fvYzqdAsBggZVlGbIs4wYN5k0R27Z16/W6OD8/P12tVs/qun7ivT+NMZ4bYy611svJZFIopcoQQuO9d6enp2G9XscvvviCTk5O3vVnYO4QLIAwzEfAZrMBAFhryXsPKSX1l+0JD239pElrfePSnwDxophh3gP2xSjamfjg7yjzExHoRBABAsWAIAk6CvggurwPAOQc0LZAXUMYC9gNyFqIraWT2GZ/qGgAYxC2Ex99JkhvFUWgD1oI2e207IoP3eP9v4FSaig8VFUF7/0gfhhj4L3HaDQabCj4+8u8Dr01llJq6NZ1zqGua1hrEUIYClm7Fijbc8Eb1iYvCkvfLbSxSMIwDPP22d337ltd7V5uCznvfybLMuR5jvl8jqOjIxweHmI+n994391pQYZ5HagjOOf6zI9lURTnV1dXT9fr9RPn3FMp5TNjzHmappcxxhURbdI0rdbrtf/000/9d999F/74xz8S534wbxoWQBjmjjOdTimEQEmSRKVUNMaEEEJQSvnttQsheKWUA+CIqPXeN3VdV1vrLKG1lkQkeNH7ccMh6O+WvfCd5/8fu99L/o4yP4WtoCbQuVZJIsgYIRAghYBEgHcOUArCGKCugSQByhLCWggpAaUg+8U5AJICSghEKSAhEQmg3fXMByqC7Bci+o/Q5S0M/4oACN4T2rZFWZa4uLgYwqt7n+2+85JhXodeyOg93JumgXMOeZ4jhACtNdq2RVVVKIoCbdsOwkifD9LbYu2Hoe8f91+WH8IwDMO8WV4Wbr4vfPS2V734EUJnxamUQpIkmEwmODw8xOHhIRaLBSaTCUajEe/PmTcKEZH33ldVVW82m/V6vb5aLpfnm83mtCzLU+/92Wg0OldKXXrvV5PJZK21rqy1rdY6fPfdd/HRo0fx0aNHPP3BvHF4tcUwdxe6urqi2WxGWZZFrXWUUgYhhFdKOSJqlVJNjLFRStXbbBDlvRfL5RJN01BZluHw8JC01kprrbgbhGHeB7riqsC2QIXnoki/UOLFDPMmEESQ6ILRVYiIAGQQIOdATQPorQhiLKLSUBAQUkECgBBQACD7EHSFqACAANEJIdgRDT5EEQTAUEDuvnti+Bj7nfV91/3V1RWqqsJ6vYZzDkmSwFr7bv545k4hpUSapjg4OECSJPDeD97uRVHg4uICTdMMAkm/7fZBuPtB6T0/FPu4GYJhGOZtcNv5fB9sDuDG1EcvevSTH/2lnzw9Pj7GL3/5SxwdHWE8HiNJEl4vMG8cIopN07jVarW+uLi4XK1WZ2VZnjrnTqWUp2maniVJcp4kyZXWehVCKBeLRf3nP//ZPXr0KD58+JAnP5ifDRZAGOYO8+TJE/rbv/3bCCAQkYsxttba2jlXCiEMAKuUktuukdY51xBRXdd15b2vhBBVmqb1eDx2UsrMGGOISBCR7K+llEJKKbcCiRRCsErCMG+BvuDa1aHEDwrItHdhmFehn1/QIBgixBgQQYgQIOkhnYNoW1BVgbQBKdWFnku53RQJIkZI0dlfSQBaSgSIYZppWMJ/wLkgved2V0S4aRHU20kIIW7YYTVNgxgjrLUYj8cgIozHYxhj2A6LeW2klDDGDIWtviNYCAFjDGKM2Gw2kFKiaZphamS3azjGODy+PwHCogfDMMzb4WX72/68Y1/4AJ4fB/r3cM4hTVMsFgscHBzg4OAAi8UCWmvO+WDeGF3WeaQQgm/btinLsiiK4rIoirPVanXatu0pgDMp5YWU8kprvUzTdG2MKQE0z549848ePQosfDA/NyyAMMwd5uHDh3R9fR2n06mLMSoikmmaiq2XFSmlIhE5pVQdYxxLKcfe+1EIIWvbdqyUytfr9XQ0GhUxxpFSKgkhaCJS3ntDREprbZIkMePxOLXWGq01CyAM8zYYks+7jIVINFgPdY+/k7+KuSNIAAoESwRCBGgrpomI4D2k80DTAEp14ocQ3YSIEJ2tVQiQRIAACAIKBKFU5621fS8BgUgEEtuu8nf7kV+b/W75fYug5xMiQNu2g2BycXEBY8xghzWdTpGm6VC8YJhXpfdvT5LkB8/FGNG2Lcbj8SCAxBjRNM1gjdX7xb8oG2RfDNm3zGIYhmFen9usCPef3536cM4NVlfGGGRZhslkMuSL9QLIdDrF8fEx5vM5RqPRu/hozB0mxkjee1eWZVWW5booisvlcnlaFMWzzWbzlIieKqXOkiS5SNP0KsuyVZIkmyRJ6qqq3O9///vw29/+9kNdBjAfECyAMMwd5vPPP4+PHz8Ozjn34MEDLJfLqJTybdt6KWUDoBZCbIQQKyFEppQaEdEIQKaUGhPRuCzL/Pz8fGKMGQNIQwg2hJB479MQgk2SZDSZTEb379+XSimp2cj8o4AtMN4hg+cVulDpPQj0ITbSM+8ZAoACkIAgCJAigkiAKAIxAsEDrgU1GqQ0guiK/ARAxAjErhuxn+xQWgIhQEnZqSvoJkAIndUW3cGN9jYRxBgzFCuur6/hvcdms0HTNNBawxjDAgjzxrHWYj6fD3kgfQh6VVVYrVbw3t8QQF4UfP6iDBAWQhiGYV6f3dwl4OY+dfc1AG5MffQ2V845aK2RZRk++eQTLBYLZFkGIoLWGtZazGYzttxkfhaIKDRN0y6Xy9XV1dXFcrk8bZrmaYzxmTHmVAhxJqW8MMZcSykL733Ztm2zXC792dlZ/OKLLzjvg3krcKGSYe4wQgicnJzEf/mXfwlJkiDPc2rbNkgpg/feWWtbIqpCCKWUMlVKpVLKzHufARgR0cg5NyqKYkxEIyJKQwhpCCF1zmXe+yzP83GMMZ9Op63WeiSESIlIABBbm6zh9vZaCiF6sWTrmsWrZYb5sdwQnkQneHQLp53X7DzPMK9DL4AMcxkEeEREEhAxIoYA8h7UNohyCPMY7K4EuskOSAFhNKAVlDadRdbWYscLdK+BRMROZ/kHfEjYD4/e7ZTfDZvuO+/7LIbeuqjvyjfGQCl1oxOfYV6XvjCmtR46h4UQ2Gw2UEphvV4PmSEAbrzmRZkg+7f377MYwjAM82L2xeX+sf3r2zI/euGjty201iLPcywWCxwdHeHg4ACTyWT4HUopWGvBfYrMm2LH9io0TVNtNpv1arW6vL6+Plsul09jjM+EEM+MMWdCiAtr7bUQYq2UKrXWTYzRPXr0yH/55Zec+cG8NXgPyDB3G/riiy8AIDx+/Jju3bsXq6oKRBQWi4UjokZKWccYK611QkSJECKVUqZElHnvM+dcWlVV1gse6KZAMudcFkLIvPe5lDJfr9el1noUY0yJSMUYVW+71V+HEDQAbYzRaZqa8XhshBCKBRCGeQ3ED2+T+OFTDPNaEA0iSCe0AQkiEAUEAnwQiFIiOPc81Hz7M901deKHVoDRkMYAiYNQEkFKkJSQQoCEAO2sez5kKyzg9q7N3a753nObiG7YYRljkKbpkBeS5znSNGUBhHkj9NZY+92//fa4Xq8HD/myLG9MifTb4G42SH//RdMgLH4wDMO8nJdNefTZTP3tXgTpH9+d+ujPHw4ODnB4eIjFYoHFYoE8z9/yJ2I+Jrbih6vrutlsNqvVarUsiuJ8tVqdrlarZ1rrZ1mWnWqtL4QQ10KIFYANEdVlWbaHh4ceQDw5OYl/6XcxzJuCBRCGueMIIYiI8Ic//CE+fPiQfv3rX9NsNovL5TLUde2JyBGRE0LUW0srG0KwRJQopRIACRGlMcZUCJFsn0uNMalSKgWQNU0zuri4yDebTWatTUMIxntvvfeWiEwIwYQQrPc+EUKkeZ5nh4eHYynleDweSy7wMMyPY3C/Irp5YZifkT4MPaVuVkMTUEeB1rsuFwTddtlviWErgEiBbuJDa0jdiSBRCEghASVBSgJSDe8RgWH64y5t1ftTIVJKKKUGO6wY42BDVJYl7t27hwcPHkApxd2azM+KMQZ5nuMXv/gFsizDaDTCkydPUFUVyrIcppD66/72i0SQfasshmEY5ia35XzsChwxxhs5H73lVS9+7Fpf5XmO6XSKX/ziFzg6OsLx8TGm0ylbaTI/OzHGUNd1c3l5eX11dXV+fX19UVXVU+fcU2PMU631qVLqTEp5LaUsrLXrEEKllGq++eYbf//+/fjZZ5/xiQLzVuFVFcN8BGzHCmlrQ0WPHz+myWQSP/nkk/Bf//VfQSkVJpOJMsa0dV2bLMu0994KIUwIwUoprbXWeu+tlNIASIQQiRDCElFa13V6dXWVGWNSIUQaY7QhhNR7n8QYkxBCsp0aGWmtR1VVTbTWIc9zobWORGSVUlIIIXkahGFeztfDCQQAACAASURBVG1FJbFz3T87FJWFQBASQYhBQBlEFIb5EezaYQmKkARQDOi3poguAB1dXDpAEUIKkJKQWkMnCYS1kGkCoToLrGg0CLp7VymArRDeb7d3hf0Oz76Lfv/5uq7RNM0wJTIajYbXaq1vdOIzzJuiD0yfzWbD9laWJaqqQghh2PZ27dy894Mg0tuv9EW82yafduHJEIZhPjZuO2+/zepqN+C8b47orwEMVle7r5lMJpjP57h3794gfrDVFfNzQR0xhBDruq7Lstwsl8vry8vL8+VyeRpjPI0xnimlzqWUF1rrK2PMSilVhhCqNE1b55y/vLwM//7v/x7Z+op52/CekWE+InaEEAKAr776Sh4fH4eqqoJSSjZNo4QQrVJKjcdjVZalqapKSyl1CMEQkVZKaSGEiTEa770FYInIXl1dpUSUEFECICWiLMaYxhjTEEIWYxyHEHIp5SSE0I5GozCdTiGlDKPRKCZJkmitOQ+EYX4EQnSeRAJ7osbNF3Xih5TwUkJKBRUjFEW2yGJejR07LCG6kPMIAUIXmOwh4IkQhgX8NjtAyc76Kk0gEgNRWkilIJTqrK8gAClAUN3PiU5IEfjws0B6bgs27YvG/eN9KHoIAUVRwBgzhJcCwHg8RpIkLIAwb5xda6x+2yyKAm3bwlo7bKfOOTRNg6ZpbhTjdrfJF4Wl7xf69l/LMAzzMbKf89ELIL3o4b0fbvdTo32WU/8z0+kUR0dHODw8xGw2Y9sr5mclxhi996GqKldVVbnquFqtVudFUZxaa0+VUmfW2gsAVzHGpVKq0Fo3bdu2q9XKZ1kWTk5OwsnJCYsfzFuHBRCG+Qjp1XYiGmpNX3/9tZzNZuH09FRaa+VyuZRZljVaa1kUhUrTVGqt+1wPJaXUZVmaGKMhIpPnuQ0hJFpru80KybbWWRkRjZqmmXjvJwBKIURVlmX97NmzxjlXz+fz2XQ6nckt7/LfhmHea/qCUV9Iul35AABECEBINFKBtEX0ARYeIhJEn9XAMK+IACBBsBQhIiDhUQOI2+mPiK0lllJAXYMGAcRCJQmENRDGgKTsJj+C7MQUpUBiRzDA3RBB9kOh+8f6rvn+fl98JiJsNpvBhqhtW3zyySeQUnJHJ/OzYozBeDzGgwcPMB6Ph4mkEAI2mw3Ozs5wdXU1TIf000nAze28P417WVg6wzDMx8L+/m9fDO5F5dtsrpxzALr982w2wyeffII8z6G1RowRaZoiz3NMJpMfZDwxzJsmhBCrqnIXFxfr5XK5LIrisizL8xjjubX2XCl1YYy5sNZeeu+XUsqiqqpyPp+75XIZvvnmm92lAsO8dXglxTAfMbvWWJ999ln88ssvxcOHD8WjR4/w+PFjobUWZ2dnIs9z8ezZMzEej8VsNpN1XUvnnNJaq/F4rIQQOoRgjTF2e52EEDIhRNq2bRZCGLVtm9d1PQ0hTIQQ681ms44xbmKMGyllkyQJSSnzGKMlIrG1w5JsjcUwNxE7N27VP4YnuwkQLxWgFKA1JEXoGKH4vJN5TYZJEIqQIIhIIAIiESJFROrWNSS7CRDSGkgTwFogsRBGQyoFCUANIej9Rd7MAOm7x+/I7n+/ILw/CQJ0xZCqqtA0Ddq2BRHBGDO8hu2wmJ+L3npNa43pdArvtxNe3uP6+hohBLRtO7xeaw2l1I3uZQA3bLF2t9N9z/v96RA+zWMY5kPntkm43ef66/1LP+nR7zf7vKVeZJ5MJjg8PMQvf/lLzGazQezobbGSJIFS6i1/WuZjIMZIRBRjjLGqqmaz2ZRXHRer1eqMiE5jjKfW2lMhxLm19jLLsuu2bVd5nm++//77Zr1eh2+++Ya2Ux+8CGXeGSyAMAwzTITgRx6QiEhi2wj8P//zP2q1Wqk8z3WWZWa1WtmmaRLvfSqlTJqmSeu6zpqm2Ugpy6ZpNs65sqqqTV3XJYA6TVM3Go1ARK1SKg0haKWUUUrZNE3NtvjDZ3UMcyti79LRF5DDNl9BSgmzLTTzqSfz2uzYYUkAoIgoBUJ8/hIvAGoloDVE2wBNA9QVUNnusT5XQEkoJUFSIgogSjHk1kgpEbfix13aXHcLIrtTIP3tPti0t8TazQMBOjus3pqIYd4ku3ZYu7RtCyklyrJE0zRDQc4YAyJC27ao6xohhOF9Yox/MRPkttcANyelGIZh3mf293G33d593X7Wx27IeT8dmiTJ0PgQQoCUEtPpFIeHhzg8PMRiseBpD+atQUSxbdvQNI0ry7JcrVar6+vrq+vr64uiKM6stWdJkpwnSXIphLgyxqzSNF1Pp9Py22+/bT7//HPHWR/M+wILIAzDvA79QSz+v//3//DnP/+Z1us1YowUQohSyhBC8DHGJsZYxxirEEJFRKUQYg2gEELkQoiVc64oimKtlNpYa+dElLdtmyVJMppOp/l8Ps+FEKm1lgUQhnkNaOfCMG+a3g4LAFTcDmsEgRgDRPAQ3oOaGlQbxNJAKPVcAJECQsrnEyAyArITRAidwEK4W7Pyt4WhAs+LJb3VVV8g2Ww2+P7771HXNcqyxP379zGbzWCMeZt/NvMRI6XEaDTCvXv3kCQJmqYB0G2zdV3j+voa5+fncM7dyAfppzx2J5z65/rX9e/TX+/mhrAQwjDM+8rLxN2X3d61u+qFjz7ro9/XHhwcYD6fYzweD0JxmqaYz+fIsowbIJi3SgghlGVZX19fb1ar1XVRFFdVVfVTH8+01mdSygsiugKwArBRStUXFxf++Pg48jGceZ9gAYRhmFdGCEE7J3Txr//6r+mbb76hs7Oz2DRNnEwmgYh8jFFXVdUAqIioUkqV3vu11roAMCaiwjm33mw267Zt1wAWIYRp27aT6XQ6dc75JEmE1pq2nQOi+/VCSClFzzv6Z2CY95a7Uixm3m+6PBDAUByyQWIUiKLzrybvIJsGwmhAa8Bo0FYAEUpDSYkgJJQQW+Hj+QSIkvKG8NELIXeBfbuf/eIwEQ1WFnVdwzkH5xy898iyDMaYwQpLKcUFYuZnRSmFJEmwWCwwHo8HaywiQlEUEEJgs9kghADn3DBJ0tMX/XYtsICbggeAoTB423eDLbIYhnkf2Lfw25/sAHDjuf3n98Xf3aaHJEmQZRkWiwXu37+P+Xw+7Pe01oPVFQsgzM8NPSfWdd1uNpvNxcXF9XK5vCiK4tx7/0wIcWqMOdVanwkhLkMIyyRJ1kqpMs/z5uLiwj969Ogu9TAxdwAWQBiGeS1280MAiIcPH9Ljx4/j2dlZACAnk4krikLGGFUIQXnva+99qZSybdumRDQCsHbOrVerVRFjXMUYl865Wdu287quF0IIl+e5BzBpmmZERFoIoaSUJk1Tba1Vig1PGYZh3hn9MlxSBEggQQAB8K4FSUAKAKrLA4myy6YhpSCEhABBCtEJH0JACwHa5tcIIRDwfPqDqHttb4t1V9gv6u5mffRWWH3oNNBZYPXFlTRNkaYpT4MwPytCCFhrh5D0vqAXQoAxBt57VFUFYwycc9BaD13NbdsOdm77kyAvEjR2xY7+9q5dHMMwzNtmV/jo7+8+t2/vt/v4rvjRZ3wopYZpjt7qKkkS5HmOo6MjHB0d4eDg4Af7TBaCmbdBjDF4733TNG6z2axXq9XV9fX1+dXV1flmszm11j5NkuTUGHOutb4IIVzFGFfr9boEULdt6/74xz+Gf/7nf+YDN/NewQIIwzA/iZ1pEHr06JH46quv6L//+79psVjEPM9FlmV+sVjIuq7d9fW1btu2zbKsLcuyjTG2AFohRCOlrL33jZRyo7Xuc0Kq8/Pzcr1eT7XWY+99prVOsyzLFovFaDKZpCyAMAzDvCP2LCDU1g5LRCAEAjUEGQMiCAHoBA0pAakghex0jO1aXm4zbDp9QwwCSRCdINJngQjggw9Gv62AsftYn6HQH9764klZlnj27BnatkVVVTg+PoZSigUQ5q2wa1XV09uyAMBisRhsXOq6xmq1wuXlJZqmQdM0t9pi7Vq/9V3NL5oA2YUnQhiGeRvsT3XsPr67f7pN6NgPOe+f6yc9jo6OMBqNkGXZcMxP0xSLxWLI/uL9HPMu8N6Hsiyr5XK5Lori+vLy8mKz2ZyHEM6EEGda62dKqXOt9SWA6yRJCiIq27atP/nkk7Zpmt0eJoZ5b2ABhGGYn8xesBWdnJzQkydP8PDhQ7FerwFAnJ2dSQAegHPOOaWUk1I6IUQbQmiEELXWuvHel1rrEkC5Xq9L7/1GSjkloqn3fpJl2WQ6nU6MMbDWSmPMcy+s7iSRzxQZZh/+VjBvAQUAFKFAoBBBMQLeIYDQAghKIkgJoTRICEj0voYSEAJSCKjtBAiALgtEAFF2kyZhv/vyAy4MvKibtC+y7FtcEBGapsH5+TmapkHbttBaI0kSWGuHLnkuljBvCyEEjDGYTqew1g4FPgBYr9fQWmOz2aCqqht2V7cJILs2WX9pG94tRLIQwjDMz8HuvmV3H7ObUwQ8n/bow8x79n9ml376ow81n0wmw/tqrZGm6XBcZ5i3xNDQSkTUNE27Xq/Li4uLq+vr64vr6+uztm3PY4xn1tozY8yZtfZCSnmdpmkhpdx476sYo7PW+r//+78Pv/vd71j8YN47WABhGOZNQgBwcnKyf8ATJycn8eHDh+Hq6kouFouQJIkPIXgiakMIDYA6xlgT0cY5t4kxbtq2LZ1z6xDCLIQwDyHMx+NxQ0Q+z3OxFT+QJInWWrMdFsO8DLFzYZifAYFOBFFE2+mQLhW9aVtIqUBaI26v1Tb4vMv/UIMIoqSEVKoLR5cEaAUiARKA6EWPvmj6Lj/sT+THdLbvdsT3galVVQ2vGY1GsNYC6DrxkyThaRDmrdEX66SUsNYOnc67Fm5FUYCIYIwZ8mp2RY4Y45Bvs2uT9aLCY3/9ssIkwzDM67Kf8dE/tv8aADcmPfrb/f7PWjtMcfbP9aHneZ5jsVjg4OAABwcHmEwmw3v3jQyc88G8bWKM0Xsf2rYNZVluiqJYLZfLi9VqdVaW5TMp5blS6lwpdW6tPQdwPRqNllmWVVrrum3bdrFY+M8++yzsNccyzHsDCyAMw7wNaCuKiO10CB0cHMS/+qu/CkopV9d1S0Q1gEprvVZKFd77VQihIKIVERUA1gCqEEJdVVV7eXnpicg3TePm8/loPB5nUkrFi1/mY0cAEH39mU8/mbdFP8Fwy+MyBMA5UNMiyhokVfc4xe66L2YCUFKBlIaUAtAaJLYZINv8kIidmfoPfAqk50Wh6P0kyG32WGVZ4vT0FCEElGWJo6MjzOdzaK25CMy8NYQQuK33ZDQaYTabwXuP6XSKtm2H1/cX7z2apsH19TXW6/UQrt7baL3qdsyB6QzDvC63CR/7Qec9u8IHgKFBobe3yvMcBwcHGI1G0FoPz/U/079mPp/faGRgmHfFthkhbDabZrVa1UVRXBdFcV7X9WmM8amU8pkx5lxKeZEkyYW19lwpVSRJsvbeu6qq3KNHjzyAKISIf/EXMsw7ggUQhmHeJnRycgIA4eTkJF5eXoaHDx/64+Pjtm3b+vz8vE6SxGqtN977UghROeeqNE2rtm3rGKMXQjjvvT8/Pw9t28aqqqKUElprZYzRUsrOUYXtsBhmpyhNg90Qw7x1iIAQENsWJCSiEADFrbKx7XhE1/GojQGMQVQS1AekSwHCtsjaW+kAoDtS5NwvuPT0HaC9N/huV2jbtkO+QlmWUErBWoskSW502jPMu0BrjclkMgSjhxBuPC+EQNM0WK/XiDGibdsf5ITcRi8KvsiXnydCGIZ5FfaFjxdZV+1Og+yKH/tTm0mSYDqd4v79+5jNZoO4sfv6/nidZRlPbTLvksH2KsYYm6Zx6/W6Ojs7K4qiuCzL8iyEcKq1Ps2y7HRreXUJ4MoYcy2l3DRNU08mk/D9999HdOIHt94x7zUsgDAM87bZtckiIgoAxOPHj+VisfDr9do9ePCgrarKA/B1XXshhNNaO+dcCCG0IYS2rmsXQgje+zgej8laS1sbBqO11jwNwnxs9O5W/Zmn2BaJZSToSFAxQhJ1NkIM8xYRsZsC0c4BQiIKQMQAFQnCe6gQoLyHCKGbBpESQkoo6k5U4zYtnZQERRqmQiS6aZC7wMuOV33Bty/S9DYabdsOuQt5nsNaCynlYIfF0yDMu0IpNWyD+zYy/TZZ1zW01qiqCt77YZKkL0Q6526IJ/3jfVbI7nvuPt8/vi+O7P5uhmE+Pm7bX7zI6qrfz9wWcA50+zhjDIwxNyz9JpMJFosFFosF5vP5kOWx/7v76Tm2umLeFdvtOYQQfNM0bVmWZVEUy+VyeV0UxWnbtqfW2lOt9VmapudJklwCWAohVtba0ntf/+EPf2i/+OIL+u1vf8uLS+aDgAUQhmHeJbQ9aSQAkYji119/Hdu2DcYYUkqRUio654JSyhGRF0LU3vvaOdcSUZBS+svLywAgeO9pOp2OR6NR1oejv9uPxzBvh2FDp5tRH4IIJgbY4GG8h96KIAzzNhFE0DEi8R4ahBgDZPAQ3kPUFWRdQTY1hGshlABphagUJEXI7ewHme3EhyIQRHfQEGIQ9O7yVn3bVEh/7b1HVVW4uLgY7h8cHAyv4Wgs5l3QF/detv3123XbtlBKIc/zoVDYti2KosBqtYJz7kZA+r4guG8fd5v4sW9lw6eHDPPx8KJ9wctE09uEj/4ihIAxBuPxGNPpFEmSDPuULMswn8+R5/kQZs4w7yNERCEEX5ZlVRTFetVxWdf1Rdu2T2OMT4nomZTyzFp7AWBljCmEEGWWZU1RFP7k5CRu3T0Y5oOABRCGYd4n6Ntvv42//vWvvbVWKKXQNE28uroKMcZWa91470spZaW1bmOMvq5rd3p66quq8nVdExGR7uCZYuajgYgwDB1vrwUATQQbAhLnYL17PgXyrv5Q5qNEgmC2216kCAQPuKYLP1cKUmvEcgPUFYLosj+gNCQRtJCg7UQIyS4oPUqB2G/ofdHi3X7EN86urca+3U9fBO6769u2xcXFBeq6Rl3XICJYa5Gm6bv8CAzzUrTWyLIMh4eHyPMczjkAnZ9+URQQQmCz2SCEMOSCKKV+8N3YFzNe1tm9/1q2yWKYu8nud3t3f/EiW6vd/cVuXseu+NHvi3pxdz6f4/79+5hOp4PYa4yBtRaj0YgbEJj3GiKitm1dURSbJ0+eXC6Xy4uqqs699+da6ydEdGqMeUZEl0qpKyHERmtdHh4e1iEE/9lnn92VIWzmI4IFEIZh3huEEERE8auvvsJvfvMbX1UViqKgNE2Dc65t27YRQjRKqQZAkFJG55z33nvnnCci2louSCKKSZIkO3ZYvMJl7gxEN6+HO7tdbtuQaU0RJgaYGAdbLIZ5m3T5M9RNH0UCRWzDy/12VElAhtBlfozG8NkIMLazcJMSeit8mC4HHVH0tlhdYSP223VfwLgDu/vbDlm73e59YaUvzNR1PYRIJ0kCYwyICFmWwVrLdljMe0c/JZJlGdI0HYqP3nsYY9C2LaqqgtZ6EECICCGEwRpr1xLrZbkhL3puX0hhQYRhPkz2v7u32eT1919mlbcrePTNBruWkr0AMp1OcXBwgMPDQ0ynU2jdldX6HCO2t2LeR4iI/j97b7IkuZWl93/nDgB8igiPyJFkWVFl9e8FadJCvZWs2GbclKy2Wa+gx8jQY0gbrbSp3LaZtGvyAWhaFc2ai7JuNYuZGZOPcAx3OP8FhkAg3CMzWSQzIvL+zDwcjuECCAfgwPnu+Y733llrXVEURZqmq8VicTGfz09Wq9VpWZYnUspTIcSJUupUSnmmlFo451bGmCzLsqIsS/P111/758+f37e+R4EPgCCABAKBW0VXBKnhhw8fOq21tdaaJEnscrl0cRxTnufCew9rbeMfrUajkRRCCGutn0wm4/F4PNBaExGFbjiBe8b2h7u6WkJrgyWY2xc43KsG3gN8eTzuOgadKMB5Dt5s4NMUPhmAhQRJBSEVpCCAqsLokgAlZZX10QQ5iFDpKvcnG2RbQdZtdlhNQMdai81mg9ls1gaNp9MpJpMJiKgN0AQCt4FdNlnWWnjvMZ1OYYzBZDJp64A0okhjjeWcu2KF1Ygk3cDjLlFjV42QIIIEAneHfnbXtuzJbe/bipl3X845KKWgtcZkMsFoNEIURa0AMh6PMZ1OMR6PMRgMwu9r4E7AzGyttWma5mmapqvVarZYLM43m81pnucn3vsTKeWZlPI0iqKLWvxYG2M20+m0MFWqpkUoeB64o4QrdSAQuHXUP6j+2bNn+PLLL/nVq1f+yZMn7uHDh3Y2m/nBYOCNMUIpJYUQdQyMqCxLeXp6SpvNBpvNxjnnWGutpJQq9MIJfHiE+9LAHYIZbC18WYCzDG69hlAKLCubLCJAoBY/GjssIeAAOCI4AKIjfvQDm3eRXeJHv7c7M7d2WMYYzGYzFEWBzWYD731ryREI3AWaHtdNAWFrbXs+L5dLnJ2dIU1TeO9RFAWklFcEkK6w0YzfJmrsukYEESQQuBtsO4d31QRqbK2aIuZNlkdf9GjabLLOtNY4PDzEo0ePMJlM2vYam6skSUKmR+DOwMy+KAqzWCzW5+fns9lsdp6m6WlRFCdCiJM64+MsiqKLOI7nZVmuiWgzHo/zx48fm++//9598cUX7h/+4R/u/k124IMkCCCBQOC2wi9evPCff/45f/bZZ/7hw4f06NEjV5Ylp2kKrbX03ouyLKGUojrwQ+v1GsYYBsBxHNNgMFBExHEcx7UQEoqjB+4F1HnvH9CtjzGq4LAVAkKIqv5HYxd0DwLEgXsEM+A9XF7CZRk4iuG1BkkFVqoKMBBBEsEJAUEECQKLSvTg2gqLcb+yQICrQZ6+ENLv6c7MyPO87Rnf2As1w1rrYIcVuNU09W0a+7YmYAmgzWxK07QNQjaiR/MOVMFNa+2VgGY3M2SbPc62nuMN24qqBwKBX4Zt595NNlb95fpiR2NvpZRqfw/7Ion3vi1oPp1OW6urhiZ7TTX3J4HA7cU759g558qyLDabzSpN04vFYnG2XC5PjTGvmflECHEqhDhXSp0T0dxauyKizcXFRXF4eGh++9vf2v/1v/4XB/EjcJcJAkggELjN8PHxMaN1TmGfZRkfHR3x//t//68p9OoAOO+9LcvSG2NcWZZOSumSJGGttbDWuvF4PB6NRgNd+WEFO6zAnYZ67y2dB8DGDsjUNkKQFso5SAAyiB+B2wYzvHXgsoTbZHBSQ0oFISTQBC1RZXlIIcCyygBhUPVe1/5g4FIEuSfHeb9He3c8cGmF1RRpbXrGr9drXFxcQAiBsixxcHCAvb29YIcVuPVss8ZqcM6hLEsMh0PkeX4lA4SIYK1FWZZYrVbI8xzGmCtZUzfZyu2y09l1LdlVXD0QCPx4bjqv+nZWu8TMhr6o0fxOxnGMOI4xmUzaGh/9oudJkmAymeDo6Aj7+/sYj8c/2z4HAj8XtfhhNptNY3t1sVgsTtI0fV0UxWvv/YlS6rVS6lxrfaG1nkkpV1LKVvxYr9eWiDyCvUDgjhOefgKBwF2g/bH9+7//e/fNN99Aaw1rLZdl6ZIk8dZap5TyZVl6IYQvy5IvLi5QFAWt12v38OFDljVCiCCABO4hnd5wXAkgIEIpJbzS8NYiBkDOVZkg73NTA4E+zGDv4MoSNsvghARLCUEEQaItcg4iCCkhtKyEEKXA8JBND8y6Fojr9Q696+yy5emKIN0aCE0QZz6fI89zpGmKOmOyzQIJBO4aWmvs7e1BSomyLGGtvSZs5HmO9XoNZkZRFLDWVhmQ9TWiOUeaZfrDu+oH7KojEggEflpuOq+2CR27xvXtrRrxwzmHJEkwGo3w9OlTTCYTDAaDKxkjQJVxFscxxuMxtNY/+X4GAr8E3vvW9mo+n8/m8/nrLMteOedeKaVeCyFOoig6UUrNhBBzIloKITbD4bA8ODiwf/nLX/wf//jHIH4E7gXh6ScQCNwZmmJbx8fH7unTp/joo48wHA65KAoAgPeeiIia3j6bzQZ5nkvvPZRSNBgMJBEhSRJfCyGCiELecuBOUHdw3zKisv6RuLwzrcM1lS1QXS+BpILyHgz3C295IPA2MNj7qg6IMXBFAWQ5WClAa3Dj5U8EL+sMEADkPUhKCCXBoiqSTo0VzrWT5m6zrchrM74byO0KIHmeoyxLMDO01hgOhxBCwDkHrTWklMG+I3BnaKyxtNZtL+3ueSGEwGazgdYaWZa12R+NAMLMrTVW11qrX1dnVwB2V6HlvmgShJFA4O25KZuj/3lb8fL+fM1zIFAJnlLKVsBoxJC9vT1Mp1McHh7i4OAAw+HwWlvNdSN0GgjcNZjZM7P33tuiKPIsy9br9fp8uVyeLpfLV9baV0T0qhY+zrXWF1EULay1q729vfTi4qL4/vvv7bffftu4cQTxI3AvCFfyQCBw1+Dj42NmZv7qq6/49PSUAZDWGs45IiKqH255s9mQtVYRESVJQkmSSADsvR8PBoO4tsMKkZ/A3YEBAtW6RxXg5coEqLoz7T68AWgrhFBVM8EBCLkfgVsJo80C8WUJJxU4zyGkhJeyFjMADwZLAd/4dScxoDTAGqRUJYR0gqIAKmss7++NGLJLCGkCvI0Ywswoy7IN9EZR1NYD8d63dh5BAAncFRprrDiOd87TePpnWQbvPeI4hhAC3nsYY5CmKay1MMbAe38lM6RrpdW3zWrOqW2F1YPwEQi8G9uE/F3CR1/w6Bcz3zW+qSfUZHtorUFEcM5hPB5jOp3i4OAA+/v7GAwGP/s+BwK/FMzsnXOmKIosTdPlarVarNfr18vl8mS9Xr9USr3SWp/EcXxeW14toihaEdFmMpnk/+f//B97fHzs37ymQOBuEQSQQCBwJyEiPj4+9n/4wx/sX/7yl7IoCqGUEnEcMwBnrXV1rx0yxrjZbGbL4F8aogAAIABJREFUsjSbzaY4OjoyDx48mIqKcB38EdwXb/27DtdWVp79pazR7R1XB5UdMzyH7juB2wuDawHEw3sHby1cWYCkAAQB7MHsK4GEGTAGXBTAcAAaDgHvQXElEEopKrGkUxMEQtwrEQTYXg+kG6Btgj+N5cdisWgDwA8fPmytP4K1R+A+oZTCaDTC48ePsbe3h7Is29ogy+USP/zwA9brNbIsg3Ou7SHezRRpXt3i6s1wwy5bukAgsJ2uULhN/NiWydh/9Wt6dO2tutOYGVJKTCYTjMdjfPzxx62VFTMjjmMMh0OMx+OQ3RG4dzjnXFEU2Xw+P5/NZqfL5fI0TdMT7/1JFEWvAJwrpc6FEHMAKyJKhRB5WZbm5OTEP3/+nI+Pj9/3bgQCPznhah8IBO4sz58/5xcvXvg0Ta3WugRAQghmZq57CApjjAKA9XrNaZr6OqWZ4jiOAIjhcCiklIKIhBAiPMUG7gRdq6tGBGHmy/F8mQzSjHMEWBAsqCokjTY/5ErmSCDwvqiO20oEcdaATWVrBSHABPhGIGEGO1vVs/EeAnVARQhIIeAFAVzlRTWGb9QUS79nIkg/aNQPxkop28BRURStHZaUEoPBoJ1fKRXssAL3AikloijC3t4ehsNhK3KUZQkpJdI0RZqmrTDYFz36hZCbnuTNedYdBm6uM7StwHr3cxBPAveZbVke/Wnb7K26WR19YaP7mYggpWwFjG69D2ZuxdCDgwM8ePAA+/v7iOMYtTVyWxNLylAaMnD36dpelWWZZlm2WK1WZ7PZ7NVyuXxtrT1h5lOt9Qkzz5h5QUQr733qnMuKoiidc/b09JQb2/FA4L4RBJBAIHBnqX+c/T/90z/Zf/mXf8FkMmHnnB+NRq4oCs6yTERRpMqyRFmWbIzxQggppdRxHA+cc9I5J4fDoY6iCADCHXDgzsBAa33VvDfCR9PrvXv3agEYIpRUBYc1GKpeNhB47zAAqg7gqlCpBVsDR4AnVPVBnIOvAxvsLMh7SDCUrHtwSwk0QXyqrN8A1NZvaAup8z2qDdINyvYDrE2PdSklnHMwxrQBX601kiRplxkOh4iiKAgggTtP17e/S2MH12R/KKVgjGmFv0bYsNYiz3NkWQZrbdumlBLe+1ZU3BbY7fds77JLDAlCSOA+8yYRsDvcFz762R3dQuZde6s4jtvMjq4FllIKk8kE0+kU0+kU+/v7qJ/3AoF7R217VRZFkWVZtqhrfpys1+uXy+XylZTyNI7jMyHEudZ6KYRYSSk3zJxLKYssy8xgMHD/5b/8l2B9Fbi3BAEkEAjcdfjrr7/2v/vd72yWZZwkiTfGeAAkpZTMrKIogveemZmNMXo+n2trbTydTuno6Eg8ePBgJIQgGboAvTXbvHoD748rGSH1q7H/afI8LBFyqnrBWzAGHqDaOiuEXgK3g8bmou7l6Swcquylysat7gVaCyCCASUIJFX9qnqCspQQUlbZH401VJ1BgnrcfRRBto0HcK13q3MOq9UKP/zwAzabDcqyxKNHj7C3txfssAL3FiEEhsMhHj16hCRJkOd5W0S9+1qtVpjP53j58iWKokBRFFBKtSJI8+raY/Wtsbrv3eHueborMBzEkMBdpFt0fJuo181S3FXUvJ/p0QgedW3HdpxzDlEUYTAY4OjoCA8ePMB4PL6SldWIlUmStDU+gsAfuM/UBc+z5XJ5ul6vT5fL5elms3nlvX+ltT6Joug0iqKLKIpmRJRqrTebzaaI47hsxI+vv/7aIzgmB+4xQQAJBAJ3nuPjY8/M/OLFC57NZn46nfqHDx/yxcUFFUVBROSjKPJSSmeMUYvFQi2XyzjLMmmtVVUt9KpvsJRSCCEo2GEFbivc/OGmVzvVhc0rwaO5c2UiMBFABEfVPEwCLKqaIIIAAQYxQxAFO6zAe4arY7QjgjhrYJlhwXDew3lX22NZwFkIZkAQpNKQWoO0BkUlSMpKBCHUFlqEpjsbU2f4fe3qz8QuG6xugLaZVhQFjDEwxoCI2uyPxlIk2GEF7htNMHQ6nWI8Hrc2Od2i5kIIXFxcQEqJ9Xrd9ibvCh/NudEVQbrB221ixps6jPQttfrTAoHbwk1iOxG1ouKuIufbsj6a8c3vD4ArIkiTxdh9DYdD7O3t4cGDB/joo49weHjYttn9LZRSQmuNOI6D1VXg3tHYXjGzK4oizfN8tlwuX87n85e17dUpEb1WSp3HcXyeJMlcKbUUQuRxHBeLxcL86le/sn/+85/d73//e/8P//AP9+3WOBC4QhBAAoHAvaC2w3LM7AH4Fy9eAFWND9psNm0gpyzLOM/zpCiKsXMullImg8FAE5FkZjEajZTWWgYBJHAb6d+VUpO7QQSmS9GDhaiCvK0IcjnNkwCIoQiQzCDyUMxtTZBA4H1SaXuXvUEdW1jv4byv3p0DewdmD0kEoTVUksAnCTiOwXEEqTWgNcB10L89T6oskOY4v09ZIMB24aMb2G3GWWvbHrUAoLXGcDhs5wl2WIH7CBFBa/3GLCcigjEGq9UKQggkSdLa7TTCRz/zwznXiord+gRd+uP64kszrmnzTdZYIWsk8HPxJpFjl5VVf3w3w6ovfjTTu9kafaGin/XRHR4Ohzg8PMTR0RGOjo5aASQQ+JBgZm+tNcaYvCiKRZqmZ6vV6uV6vf7rfD5/rZQ611qfjcfjWZIksyRJVtbadH9/v4yiyKxWK/fZZ5/5zz//PNheBT4IggASCATuFUTEzOx/85vf2PPz80JKSWVZElD5PwNIpJSDKIrGzrl4sVgkAESapnx0dMRPnjwZTCYTUkqFyE/gVnKlvked4YE2w6Mu9FwPt+OoLtpKAgSGJYFCMAgSngkxPKJghxV4j3TDIk0tGw/Agy+DHgAsMzzqYuiCICINnQ3AgwE4joEkBukIUApCVgXUUWeKXGZN1e/3zAqry7Ze5M2r6bne1DLYbDZ4/fo18jzHZrPB48ePgx1W4IMljmNMp1MwMx48eNBmSfVtr5qXMQZ5nuPi4gKr1QpZlgHYHkTuB4p3BYWbYHOTgbLNVqv7eVf2VyDwLvSPo22ftwl5zTzbatt0j/H+cLeoudYa4/EYDx48wHA4hFKqzdLaZo8VRRFGoxEODw+RJMnP/J8JBG4nzjlbFMV6uVzO1+v1yXq9fpnn+ffM/EMURSdRFM2UUrM4jpfMvLbWplEU5f/6r//qBoOB++KLL4LlVeCDIggggUDg3lGLIO6bb74pAfByuQQAWGuJiAZKqQERTbz3yXq9TtI0FXmek3NO7O3tqeFwKBGuj4HbCDVFzusHyM6kruVVJYTINuOD26CNhyMCCYLwAhBVRJg8Q6G2LHg/exb4EGmCKqiOX0dU1a5p6tdwdaR7ZjjUgggzHFcZIawkVFHAZRlslkHGMXSRgJUGqaomiKCqIDr72ijuUgupa4LUJ9U9Cxxu66XbzQbpTi+KAhcXFyjLEtZaDAaDtrd7d5nuKxC4r0RRhMlkAq1129u8a3XVL3ReFAXSNIW1FsYYlGXZLgdcnnc3FYNu5utP7wae++f0thojXYIoEngT22yqmvHdefrvb8oA2XbMd5ftvoDKYm4wGGB/f7+tR9UUK+/P26010hRBD2J94J7D9TnATU1TAExEvizLTZZli/l8frJcLn9YrVZ/ZeYfiOjVcDg8JaLlYDBYjkajtVIqK8uyWK1W5e9//3tftwEEASTwARECfIFA4F5CRL6+Sebz83M6Pz+nNE2FUmrhnEuklMM8z3VZljrPcwIg4jhWxpjEORe9580PBK5BTbf1JlhLl0IIcJkJ4ussEN8MS3FpfdX0hvcARG234RmKRFVg+v3tXuADpKpZUx2nRghYIeCEAIuOMAJciiHe16JIdeS7soTLC5gsg9pkUFEMozVAVZCeAcAzKNKAIJAQEETwqAKYoq6bg7r2yH1jV/2BbiC3KTCbZRmstfDeYzQagZmR53krfiilMBgMkCRJG5gKBO4jSilIKTEcDt+qdkee54iiCEVRtOdQmqbI87z9vKswdDezozutER+78/Tr+PTb2db7vkuwzPqw2fb9CyGu1OzYNn9fgOhmJe0SNLZlhXTnadaplEIURRgOhzg4OMDh4SEODw+xv7+POI7fSsTrnzuBwH2DmeGc88YYl+e59d5bIjIArLV2sVqtTubz+V/n8/kPaZr+NYqil0mSnIxGowspZaq1Tr332WQyKT799FNDRO5971Mg8L4IAkggELjPMAD/ww8/uNFoZIQQhVIqFUIsnXMDKaWWUmohhFRKaa11IoTYJ6Lggxm4dVR91RkkCPB8aeFTZ3SwILAUleDRvtdZIEKARPWQ6EUV9vUs4Go7Ic9cF1K/f0HgwO2FUWV9FFKhEAKFFLBUiXeNURVxHeBAx56N66nOwRkDV5YwWVbV/pASHgQJQHgPOAtyCUgrkBRVZggRZB1gbLJK7jPdINS2YFHTu917jzzPcXp6ijRNEUURnHNQSmE4HOLhw4eYTqfQWoeAU+Bes8tyahvN+XF4eNieS845rNfrNjOke9517bOaV7emyK5x/Vo+23rv3yTY7BJEd43btXzg9rDre9slkjXL7BI7GrqiSN+Cqvu5WXabVVV/XX2hRAiB4XCI/f19PHnypK3j0dhfhUzDQKCCmWGMcavVqpjP51me5xvv/UZrnTLzLM/zkyzLXjnnXjnnXgM4J6KllDJl5ixJkuLBgwfm6dOnDuFBL/CBEwSQQCBwb6mtsFCWpZNS2iRJSiLKyrJcaa0ja62qhQ+llIqVUkMAuffeOOccdXjf+xIIAFd7xHtcBi4byytICVIKkNUwVCWGsBSAE4CSYFdbDHHTm76yBwIRwEEECfxyMKHN/iilhFGqEj+IQCAQMwQAiTppiah9MWofK+fhjYHNcxRKgUUlgCgA0nuQcxDOV7VBoggEQCjVttdkVPnWDet+H//beuY2PXGJCGVZYjabYbFYAKiK0DaWQEopxHGMKIquWGQFAh8yQghEUYSDg4O2rs56vYYQAsaYrQJIV9zonke7rH6a+iP95Ru2ZXx0x98U8N6VlbJt/ncJuAd+Gt70P78p06d/ve8fJ9uyOZrluoJGv/5GXxDprq+xfuuLJM1w8y6lhJQS4/EYjx49woMHDzAej5EkSVsEPRD4gGltr5xzPs9zs1qtstPT0+VisVhYaxdRFM2J6BzAiTHmxFp7prU+AzAXQqycc5ujo6MCgEnTtHGSvd83uYHAGwgCSCAQuNcQER8fH/Ovf/1rt1qtzHQ6zbXWaVEUSkqpmDmqxY8BM4/yPF9tNpuEiHQcx0prrWS4Ew/cEiqnVq4dr+hSCBFVxgcpCVYK0ApQCqQ0SFuQdZUVEBFAHmishNiDyQHsAE8ISSCB90XbG1pKUB3ck1wVQRdciSBNbRCubd4aSzdvLHxp4IsSVmXVuSCqlyQBFgJCSqAONlanUJX9gbYndXVqtVXS7yn9XuBNMBVAG9zK8xzOubb4vNYa1lqMRiNEUQQpZWuFFbJBAh86UsorIkVZltjf38dqtYL3HsaYK5kbXfuhZlnRXpuqAHL3HGxEFSJq528+d1/bevYD2wtXbxNcdrXRdrR4g4VW365olygTuMqu/2v3O+6P686/7fvqf25Eh+76uuJYV6gAsDXbo3k1x2Vj7dbU4WiOzWYagFYM6YsfTdHz6XSKw8NDTKdT7O3tYTAYXPlNCgQ+VBrbK2utzbLMrFardLlcLmez2XyxWJyXZXmhlDpXSp0ppU6J6EwIMSOiuVJqCSAlohyAiaLI/Pa3v7Woan6Ep7zAB00QQAKBwIeAL8vSxXFshRC5UoqUUmytpaIolPc+8t7HWZYlJycno7IsaTKZYDqdjkaj0TAIIIFbQxNY8L5K1iDU9leiChwrDWgNEUXgOILwDvAOxLVllpMQrvpMzCDvQdZUgoizgA+2sIFfDmJAgBH5SoAjloCQ8FpX9m1c1/voPK5Vh32dBdIEDwEQe3hTgksFVhqsCrCSYCkhlWqLokPVQR2qhUO+LLQO1IlQ7+Of8TOzyx6nGzyVUl4JXjXBr6ZGyNnZGbz3KIoCDx4c4eBg2gbAAoEPmUacaLKlnjx5Aq01Hj16dKUYevO+ywKrLEukaYrT01Os12sYY9pzsglkdwWTbW126/t0p3eFkDdlunXttprP3X3dtv/bPvdFlSCIVHSFjK64tMuqcJvlWf876dfy6Nfs6C/Xz9zofk9dwaMrgDjnrrySJMFgMMDDhw/b7I3+70e/7eZdSonRaITDw0OMx2PEcRwyPwKBGmZmY4xdr9f5bDZbL5fL5WKxmOV5fuGcO2XmM2Y+d86dAziL4/giiqIFEa2SJElXq1VRFEW5Wq3cYDBwv/3tb9uSeoHAh0x4Ygncdn7SO+X7YG2x5eHh7u/Uz8zx8TE/e/bMf/755/Y3v/kNAUCSJFwUhSzLMlZKDay1g+VymRRFMVqv1+ro6EhqrUWSJBGAUPE18N658vBLlW0V1T3hSQqISIO1gogjwBrAxpXNlXeXpdKdh/AO5PylACIIgj3YmarIdAhQBH4hCIAEIaoFOUEAKwkfRfBKXRY/56pCTSWYVMsJACwqwYSotstiBhsLGANYCxgLMhZkLYT3rfDXFTwYgENlh+XZ3+sf1G3ZH326gdVur3RjDBaLOcqyQFkWICJofdUKKwQ3Ax86TfH0hw8fYjKZwFp7LcNiWyZGc/6s12ucn5+3RdTzPG8D201weFuwvHlv5m1El+70RtDYljGwra1+BsJNGR39wHw/y6C/3g9JENn2/95lX9Udt0vs6I/rC1p9G6vmuOiLX9u+I2C7YNIVQ7rfr1KqFfyOjo4wHo+vLLdNcOuuT2vdiihB/AgEKtsrAOy9d0VRlIvFIn39+vV8sVhcZFl2bow511qfaK3PiOhCSnkhpTwfjUZzrfVaCJEul8vCGGNPTk7sdDr1v//9733I/AgEKoIAcn/YdgdJx8fHV0b8+c9//pvvNJ89e/a3NvFWbX711VfvtK3ffffdG+f/5ptv3qXJW8U333yDv/u7v+N/+qd/wtdff31l2meffXbtR+3Fixf4/PPP2/HPnz/n3o32h/RDyH/605/8ixcvMB6P6ezsDEIIJiKllEqEEANjzCDP82Sz2YwARFEUJcaYkfd+/MbWA4FfAiL4+sFR1J8ZVfFzUgqkNRBFVYaH9xC+Km4uQPBUFX+GMe00yQzlPYSpesazIHhj4Lh5+KVf3Alo2/p+0gvV2+7Qh3R1/KXpfAfNv1mAIJWE1xHUcAgVJ2CtIbiyvxLs4QAoBgwzJFeiBRNV9W2EhBASgkRV3BxoBT7ROd6pCcIQgaiazxNBgOH9h/Olbwto9gOf3WDUpS1PAWtdXbx2hCRJIITAYDC4UhckEPhQaeqBNAWe32Q/1YWIEEURiKitwaO1bq2yGoutvkjZrBeoLIeMMSiKoi1M3bTdiCPbxMp+hshN27mNbbZKzfL9OhPbbJ362/I267pNbPtf7fo/7hIuuuO2TeuO707bZW/VDHdrcnSXbz43mUvNsda02QgezXG0zQJrMpng6OgIR0dHbQ2Pbf+bXfvSHMPhtyMQaO+1nLXWFkVRrtfrdLVaLWaz2cV6vT4ty/JUa30qpTyRUl5orWdEtCCi+WAwWHrvs8PDwyzLMvt//+//dcfHx03Nj9t30QwE3hNBALnb0PHxMQGXwsazZ8/w7bffEgD88MMP9PTp03bmly9f0ueffw4AOD8/v3J3uVqt3ios9Omnn+Lbb799p4389a9//cY2v/rqq2vjT09P3zX29sb5X758+Y5N3h4++ugjnJ6eMgB89tln+P7779tpaZoyAPzrv/4rDg8P+cmTJ1wfC3j69CkDwFdffcV/+tOfGLgqjhwfH38QP4xUFUT3L168sEmSsDHGM7NSSq299wMAiXMuLstyWJblwHs/ATAlouAJFLg1tA+vqHqsc+XjUxU81xoySUBc9XRvbH68qKcXBeBcVRS6DggL5yBdDI5jcJLAedv2tm8FkL9RBXmXxW8SQH7cRYpu/LgTvjbw49Z3vcGfkb6y8P4u6zfGr1qLqU4ADKhs3JSGiGLoOAakBPkqq0OA4ZjhGBC+EkMc1wKIIHAt8AmtIZSCVApaCkgpIAVBUpUxIoiqjSOq7K+EqLKg+t8b8weRCbWtR3qXJuDaBNiMMW19gvl8BimrIs/T6RT7+/uhB28ggEsR5MfQBJYfP36MwWCAPM+viR7bhI/mPC2KAuv1uhVCuvZbXautZlx32i76gumurI5m3m29/fvZADfZcN2UHfI24sdPkVXyY0SWbUH+7nBfAHqb/0N/X3aJH9syQBoBo79cVwDp2rZNJhMkSXKtja4tYt8WazgcYjqd4uDgAMPhEIPB4B3/a4FAoMF7z9Zam6ZptlqtNouKi6IoTsuyPPHev5ZSvtJan0VRNFNKLZ1za6312hizefjwYa6UMuv12j1//tzXMZ5AINAhCCB3EGam//bf/hsBwGeffUaz2Uw8ffoUL1++pFevXtHh4SEuLi7oo48+QpqmNBqNCACePn2K5XLZ3Em1d1QPHz7Eer1+67vFwWDwTneWq9UKh4eH7ec0Ta8s/91332E6nd7YRn+ZbURRhCzLds63v7+P5XL55g2+pZRl2f6IzedzEBGGwyEDgNaai6LgX/3qV5hMJpznOQPA3//933OWZQwA//Iv/8Kj0cgDwJdffskAMJ1OfZ0lRHWGyL3+oaz3r7kh8L/61a8KpVQWx/HKex/XxdCHURSNlVIHSqkiCCCB28KVh+Q6G0QQtQWhSWuI2EHWVZwZVY0DlhKsCyDSgKmtgFzdM54Zkqth5z2YfWsxRERtYJi6dRHeIrhAW4ffInCxbb/b/b8+7q1a6W/vGza/uQry2wgIW2fpr2DLTFu24W8K2lx+OfXnn+NS3pct+nR7OG8dXbVSC3NVi9RuukdV00M2xcpJQHoPywwJwNXHqEIlfrh6i6paOJXIR0oBSkFqDaUUpJRQUkI2AUSiqmZOE7xrAlFNz+hqA+9/j4AOuwJwzfhuT/NmnDEG8/kMeZ4jy7LWC74pkB4IBH4cWmuMx2N8/PHHePjwIZxz1yyT+lkU3UyL5XKJk5MTpGmKzWYDY0w7vanx0y/I/iZLpoZ+0P5NAkU/wH9T0P9dsk128VNmhryrRddNFlVNO/0MkJuGm8/bskW2iRnd4b5NVX9cV8yQUrbFyB89eoSDg4OtGSu7hpVSGAwGGA6HP1r0CwQCLb4oCjOfz9OTk5P5fD6/yLLsvCzLUynlidb6VRRFP0gpz4ho6ZzbKKUyY0xelmXxz//8z/bbb7+1H0JMJxD4sdz/7m33Azo+PqZG7CiKQjx58kTkeS6MMUIIIWezmfDeC2YWWmtiZqGUImYWUkoCAGMMWWup+WytpSRJYK0lY0x7LDS9P7ZhraU4jmGtfadjp79Md/hNN0zOOXrbm6qbtuuu3piVZdkO+9qjQ0rJzTSlFCul2DnXvg8GA++cY601Sym9lNLnee6llF4p5ZVSPk1Tf3h46BaLhXfOudFo5B8+fOhPT0/522+/5Xv+40kA6H/+z/8Z7e/vj5h5P8/zaZqmD8qyfHJwcPDJ0dHRp7/+9a//v+l0+ul4PH6otVZKKSmlbOLD9575fI7Xr1/j3/7t3zCfz5Gm6bWHtZt6Dwd+HpqArQCq3vHOQRoLZQxUWUIUBURZgvICKHIgL8BFAbJVLQRylfBB3kPWwWXZtAUAqIQVwqUJFon6gRjUGe5sU38bt37+kZcTvvJ2JTmj3+K1ED01b4T+pDduz1tlUdA77FYvuHFNp/lbBRDqDF+34XjrprYFw3cMX53/asZQO0xb5qXLI6L5zqphgieqMpdQCx3McN7DM8MDsJ3hZpn6hxFUiyBCa8g4hogjiCSBHAxAoyFoOADiKuPJaQUrBUrvUToPy1W7zJV13IeQAdLlpl7dV3sUe3hf9QtogrWPHz/Gxx9/gvF4DKU0mBlaKyil6sK2KggjgcBb0FgONa9t91h9MaTBOYfVaoXXr1/jr3/9KxaLRfsM0RUxt7266y7LEmVZXhNfuuvetj3dz7uyF97F5qhvk7XNum/bem/atpvYJt7cNO8u8fgmUeNN6+5neADbs2q2ZXl476GUgtYacRy3tlL92h3dVxzH2NvbwyeffILHjx+3mXxv2oeuMNPYszUZg4FA4O1hZs/MzlpriqLI1+v18uXLlxevX78+n8/n5865M2Y+1VqfSClfJ0nyUms9i6JovdlsCilluV6vzWw2sy9fvmxsrwKBwA5CBsjthgDQs2fP6OnTpyJNUzkYDCSq7615V2ma6iRJpBBCOueUtVZGUSSstZKZBQDhnCMhhJBSkhCCvPdERK3wIUQV0VJKtTdQAOC9v3InQ0TUiAz9aX2aNgCgKIp2Xu89velBuNt298bPObdznW/aHmvtW897m7DWQghRhbTqf0SdItmMZ+ec994zM3sAnOe5JyLvnPNKKcfMTkpprbUuiiJrjLGj0chaa02SJFZrbYQQbr1eu/F47P7whz/4Fy9e+OPj4/sqhDAALsvSJUlijDG5lHKjlFrleT4yxizTNJ2fnZ3NnXPzPM+Tvb29wXA4TIQQItzgB94n3Qdz3wQUlKoKmNf+4ZCyeikJoSMgiUG2sr9qLLAEXxaeroIcVeKAaI5vuoxeV9kkV2WM7kXhMgR+fRr1Pr9h73aO7q+X6rSU69txXQDhrXZeP4EA0lcxdje0fWz7r6Y3/o+2hCB6E7piTKfX6FtsIfWGrgXAcfW7bYe59013Dp1m/6p5qDu5t0ZqC5KDudUdRPOZAcmVBZZnD8lVdo7zVSYJc3N8VrVAWhEk0pBxBIpiUByDogiQqsqIqg766oegH9xpToQPjJuCi0JQ+z16XwVSrXUoS4Msy7BYLKB1hNVqCSHFWrMxAAAgAElEQVSqXuZJkmA8HmN/fx+DwTAIIIHAW0BEUEpdeYZ6W5pAd1mWMMZgOBzCGNO22xUftgkg1lrkeY7ZbNYWYAeu2mx13/uCRt9Sq2/3tK2t/rL9rIluO00Nk/58u5bf9vlt2Zat0Z3WbE9XCNkmivTH72q3n7Wxbftvyu5osjoGgwEGgwEODg4wGAygtb4yH3DVNiuKIgyHQxwcHGA8HmM4HAYRIxD4BfHee2utybJsnabpcrlcnq/X67PNZnNWFMW59/48iqIzIjqTUp5baxdJkqyiKMrOz89Nmqb2008/td9++60P4kcg8GaCAHJ7IVSZHwJVHECtViv15MkT5ZyLsiyLjDGR9z7WWscAdPNSSmlrrSYiyczSOdcKIVJKcs4JIiKllGiEkEYAqW/oqJMe294FMTM1781wgxAC/XG9m7h2mpSSmnallK0/bZddAkV/fH+du7YFQPsQcNOyfys/VihotmXb8vWNLdc3/kxEXKe0N+IHSyk9EXlfdcv0AHwthljnnJVSGu+9ieO4dM4ZIUThnCu997nWulBKFcYYI6U0xhj7l7/8xQJwv/vd7/yLFy+4bhP40V24bycvX77kjz76yI5Go2Kz2WTMHHnvV5vNZlGW5Wyz2ZzNZrPJdDqNPvnkk6lSSsZxrN/3dgcCzNwGopmqXvNCKTgiQBCElBB1T3gYWxVGt/ayKHQtflQCCLUyR2N7RbgeoOBOMP3ND8iXkkg3YP4We7Zjf69Pba/g10SQbWuja4LD2wggb97NHy+AoLM9b3thvS5LoL/zvfbfNftj+/jL/1b3b2+hNvjVfAedwM211jrCSHcz68wL6sxJ7MG+yk7yTXZGPQwieM+t0EOits+SEqQVhFZgpUBxDI4jINLwSoGFqI/n+kX8IWoeO+n27q0+N18z1T2KAaUaOyyL5XKJoiggpKh6kVuHyWSChw8ftT2S72oWbiBwVyCqiqgfHBwgiiKUZXmlQHZfjOgLDFmWYblcIs9zLBYLbDYbALiSOdIs12+zL350p3ft8/rz189sW7NauuJKI7Y0Isg2caUvgvyYQP5NgkdDdxu2ZUo04kh3XF+46Nfn6I57G9GjeW+yhJqX1hpJkuDhw4eYTqdXBI1+210LrNFohDiOg/gRCPzCMLMzxuSLxWI2m81Oz8/PX2dZdmqMOSOiC6XUhZTyQko5l1LOAawHg0G22WzK8XhsZ7OZ//rrr0O9j0DgLQkCyO3imtVVHMeyKAq1Wq2iyWSil8tlRESJtTYmosR7nzDzwFobM3NUB3Aj770mIk1E0jmnAAhmFkIIwcwkpZRxHMvhcCiTJJFSStHplXNN9Gi2rzuOmal3k7tVjOi304gYu4SKXW11pt0oXryNsPFziB8N7yqCdLdl27Kdhxdu5mkyQWrhg621rigKl6apdc5Za60D4IQQ1jlnnHMlEZVEVDBzKaXMlVK5EGLjnMuKosi994W1tgRQKqXMZrMx6/Xapmnq//t//+/u5cuXDMDXGSHt9txlnj9/7v/3//7frixLE0VRsdlsciJKi6JY5Xm+WK/XszzPD8qyHAyHQ6WUUkQkazssIaWkm47VQODngLkT4qe697wgONTFTT3V9RBkFfyNHOAc4Kvi6PBVQLnJ72hC2kRVF33PuFYDZFv2xTYxpBse7/bxf7uLxQ2ZEr1YP3dH9IWaLdu1e003bBm/SSjptX/jTm6VLt6JG/477eB1/ePtLk916Ol6r9rLiXUEnHr/bupMbrI3uvM1bXbEjs7fTrP1LlyqTu221FkgQJ21VLdJ9Q7LZtvBVRYI1cXN5WVhdFYS0JX44Wvxw6ESUbpZIO3wB3xZ7wYXd88jUP23qvuToqh6nHvv4byDNRbGlJBCtgE45soySykJIUI2SCDwU9NkjwwGAyilrgTG+8IEcDWwT0TYbDYgIuzv7yNN0zZzvps9skv82CaAbBu+SSjx3rfZK9771oKrmd4t6N5dbpsYsm0du7JBuoJCVyzot9dvoy9udPexEX674k933u7nbk2Obe1uy95ohvsZIPv7+9jf38fBwQEODw8xHo+vCDP97W+2T2sdsvQCgZ8RZvbOOTbGeGZ2zOyFEM4Yk+V5vkzT9GS1Wr1ar9cvi6I4Y+ZzKeWMiOZKqblzbiWEWO3v7282m035ySefmBcvXnhc1ja983GZQOCXIAggt4MrwkfP6koTURTHcVyWZczMAynlQEo5YOaBc27ovR8yc+Kci733MYDIORcRkfbeKwCKqqdV4b0XAITWWsVxrA4PD+ODg4NoOBzKThZCG5Rvbnh3ZYL0vVz7N9d9sWJLlsi1J+w3CRw3CSdvy10UQDo3sNx/ZVlml8tl6ZwrVquVMcYYqop3WyllycwFEZVFURRCiJyZM+dcJqVMjTEbrfWGiHIiyr33hXMuHwwGBQDzySefmNls5qIosqPRyH/11VdNdsmPzni5RfC//du/+X//7/+9Wa/XhbU2I6LUObcqy3JhrZ1bay+cc4M4jrVzThZFIQ4ODuLRaBQJIWQQQAK/NN0HfmYGhKgCt0TwggEWVTzZOUDVXbfreh9cd+UmvswiqRqtQpmXckf9IF9P7harrsSPLdH2lk4AovP3TbQhaOqN7Ass3GQZXFvdG+/+r56u2+du5+GO0LKrva5AtHXWN8oWb89N285bx777Kjp/W6GNutP6w5Vo1p23kYwIbULH1Y2jy/9bI2ZUbXQaroNhXe2lOuYaM7PLYfZ1b+FKtavWLSUgqMoIUZUdHEsJLwW8EHBEVW0RAB6XIkgrfnzg6SDbAn+X505jl8d1ZkgVfDPGwjkHay2stSAiSKGgtIa1BtZa7O/vI0kGiKIQaAsEfg6aWgw/JuOqeabbbDZgZoxGIwDbxYo3vXczPN5mmUb8WK/XWCwWMMZcEzz64uy2Z87+566gsY1dGRxdUWPbPM1wd75mfxtbqclkUtdAkleWba6Z/W3alhXSbb8vlGxbZn9/Hw8fPsTh4SEmk0n7HQYCgfeLc47LsrSr1aooiqJ0zpVSyoKZV2VZzler1Q/L5fLVer1+WRc5n0VRNCeipRBiORgMNlrrzDlXLBYLs1gsuvU+Puyb1kDgHQgCyPuHjo+P6Xe/+504PT0VAJTWWjnnNIBICJEIIRLnXMLMA2YeMfOwI3wMnXMjZk6894lzLiaiyHsfMbNGXSekzvwQACQzU5IkOo7j+PDwcPzkyZPB3t7etTvlfoZHf9rWnXnDzejbCg9vMd8HE3TeEoS4UpODiHixWJRSymw+n28A5GVZlkIIR0TWe18SUUFEpZSyIKJcKbUBkAkhUqVUCmAthMiYOVNKZVLKzDmXCSFy51yplCofP34snHM2yzL31Vdf4YsvvvD1Tfmd/dElIvzpT3/y33//vYvj2AghCiFEJoTYCCFSKeXKe7/cbDbjV69e6TRN5Wq1knXBeaG1lu9S0DEQ+Km4EhCoA7aOqA0AAwAL0QodTUCXuCp67nxV+6Ntr33wvwxEdwWQtt1uoP2NGRLvdqHuijG9na1n4CuiRyOYdLbyXZIwdo68ltGyMxjeFYjesGLe0u47cn2ZG8b8yKtyv1h8I2pwIzzUqsa2ovLdjA/qfGetoNZZQ3uMdYbbze6Or8URqhWS5vtoBDgGQHwZkG+OW67PBQhR2V0JAS8FHAl4QXAgeKrstJxvAvnVTuwKlH1odAOHjU1Nd1qT1XEpHKkrx7hzDsvVEsYabDYpjCkhhIBSKthhBQK3EKUUhsMhHj9+jMlk0hZQb9j2TNgVCPoZHtvm7X9ulrfWYrVa4eTkBGmaYrPZXKlfAly9FvWts960zrcRQJrPuzI/usLIrmWbDJzJZIKPP/4Yk8mkrcPRnW/b9vTH96+5fVFk23xxHLfiS7jOBgK3B2ut32w25vT0NF0sFmmWZesoilIimgOYFUXxiplPhsPha+/9TAgxk1IupZRr51xqrS0AlN988419/vy5reMv4YY1EHhHggDyfqFnz56Jp0+fitPTUwVASikjY0zknIuttUPv/agRO4hoGMfxZDgcjrXWYynl0Dk35MoCK2HmyFobA9DMrL33mpklEUlULhGiFhbEeDzWdfbHeG9vb7i3txe/68a/jZjxc3WO/zkzOG47O7JEiqIosoODg5SZC611K4BIKQ0RlUKIUkpZCiEKpVQmhMillBshxIaZ12VZpsaY1BiTeu9TAKkQYgMgGwwGWRRFubXWjMdjI4Sw33zzjf3LX/7imdnfYRGEnz175gHgxYsX1hhTAigAZFrrtRBi5b1fWGsHs9lMFUWhpZTR4eGhrm3n7up+B+4JTezYA5BCwNcP6a7ODLFcXfyZqxoKop6XuCkyXXlZE2+xvBFXP/+iR3tn1ZdB/U46QTdbYMt2XRv1DtkZb2OZcbmZnQyQrVwqRtc6BNzY8s28KTPlx7RN/SG+no3T7EIrhnSX72oenZZacaKpLbNDsGJciiyVaHc1e+QyMYMvF2wCb1e24zIzCk2tDyI4Inigyvyg+t1fZp8wQh2QbTQ9j4moa2taT2uuKICAAMmrPbWttVivVyCiulf0uO4NfWm5EjoRBAK3gyZzZG9vD6PR6IoF1duwpdPbjYJIF2NMW7dkvV7De99acHXb39XmDgeCt972Znu7Yk53H/oZIX0RpBmvlML+/j6m0ymOjo6wv79/RQDZdX/xJoFm2/9v2/JSylZkDpZWgcD7hWvbK+ec32w2xXq9Tufz+eLi4mKRpulca73QWl8IIS4AnAohzuI4PvPeL4hoZYxZJ0myOTg4yIwx5rvvvnMAXBA/AoEfTxBA3iPHx8f09OlTMZ1OVVmWOk3TKEmS2BgzKMtyKISYeO/3AIydc+MoisZRFO3v7e3t7+3tTaIoGnrvG/FDO+eiWvRQzKy897IWQIT3XhJRU7ychsOh3tvbiyeTyWg4HA7iOA7dRO4ww+GwHI/HydHRUay1LiaTiSEiT0ROCGGFEKZ5SSmNlLKoBZGciDbW2vVqtVotl8uVMWblnFtFUbT03q+VUmsAuixLFcdxbowR1loBAL/5zW/sH//4R6CKgNzJH+LqtGAPwK1WKzsej4soijLvfUpES+fc3BgTF0WhrbXRaDQaGGOGdcH5O7nPgftFI3p49Gwl6nGeAIGmuDm34kdt2HAZPO5kgQBXD+42GNDO25nx56DX9JVMjI5F0dagwBtHXGaP3MgW0aLajGtZeTe387dswxubfKP0ciPXRI/OUJNRUY2jy2nUHW7mvb7mNuOjnadNs7i+tsuVXmn/8nvvZHk009rNq0uu1+cB1WOac4Cb8wAED4ZjXNpfMcOxD9ZXb6AfDLw6raoHUo2u3okI1laWWM5ZpGmKxWKB4fC8zRxpeiiHXsqBwO1ACAEhxLWMhV8CYwyICEVRYLPZQGvdjgOuiynbxJD+9ekm8aDLTVkX/XHAVQuq7nJEBCkl9vb2MJ1O23oc7+P/GQgE3j91zQ+bZZlZr9fpYrFYrVar2Wq1Ol8ul+dKqQut9ZnW+kJrfTEajS4Gg8EMwJqI0vV6ned5XiwWiwKA+6//9b/e2XhLIHBbCALI+6G5ExPT6VQBiLz3sZRyUJblkJnH3vs9Ipp67w+Z+YCZJwD2kySZPnjw4PDx48f74/F4SERRbZclasGjsbpq6n1Q897JmiCttYjjWI5GoyiKotD97o6jtZb7+/uxUkqUZZnURdBBRF4I4etsEC+EcAB8LYo0RdLLLMvWAOZpms6893Pv/VxKOSeihXNu4ZybSymXWZalg8FgU5ZlsV6vSSlFX375pfn888/5+PgYuKM/ykTEx8fHfm9vzzKzGQwGmbU2jeN4XpZlIoRQzKyjKIrjOJ4opQoppXvf2x0INHBtD9QNUPs66wO+Gi+o6rUomoBBqyc0RaXR2g8BvZOZr4fbf7a8rzby3Vl9dxuaYMS2rJVt3LidbxZB/rb2f7rF/lYLra1tXmlxe7CHaxsr6s56ZdnOd3Bl8PKL7AoXV9rqtdlff9XCZRYNOkJFM60R9i7FGF//rwhgqhJG6qB7JYRUnz37tknest+B7Xjvr2SCXBcEBaSk+t3BewkiwmaT4dWrV8jzHGm6wccff4z9/f0ggAQCAUgpMRgM8ODBgzYTpF8no5/xscsi6qdmW1bILrGlyaIZjUYYDAYhwy0Q+ICx1vo0TYuLi4t0UTHL8/ylEOJ0OByeSinPtNZnUsoLKeXce790zq2Gw2FeVh6EZVEUFoD74x//GMSPQOAnIAggvyx0fHxMf/7zn+nLL78UAPTZ2VkspUwADAEMrbUTa+0egAPv/RGABwCmw+FwfzQaHezv70/39/ene3t7++PxeCClVI3AgVrkaLI8AKDz+UrxcCIiKSVprYWUMtyd3XG01kRESiklmFlzRVsvpM5yaGqHNOM8AHbOGSHEZm9vb5xl2ch7Py6KYszMQ2PM0DmXOOciIUQkpYyZOQKwMcZIY4z49NNP6T/9p/9kfve73/kvvvjCN+2/3//Ij8IrpfzBwYFh5tJ7n8VxvGLmARFF1tqBUmpERGtrbZZlWRFFkalT3gXVvO+dCHzYMC6LmXvv68Bv0zO+Pjz9ZYC4zetoutS/05n7M53mO7IltvbGfJuAx98igPzMvNu/++16s77bBlyRtK68VdN3L3rTVlSCWke4eJdN6iywVaBpj9+rIkv1ueubdbnyxoLL15JJJRheTruLP1jvi12Bxsse2ALNLYAQBGYJ7ys7rOVyCV/XXBmNRq0FllIKQohg2RIIfKAQVbZ4o9EIURTBObdT/Oiy61r0Y3gXAeWm62DXhioIIIHAh4X33jOz8967oijyNE3X8/l8uVgsLlar1Zlz7jURncRxfBpF0ZmU8lwpNSOildZ6XRRFppQyAOwPP/zgptOpD+JHIPDTEQSQXw569uyZ+OGHH8R//s//WQCQdcHyoTFmBGDsvZ947/edcwfOuan3/oGU8mEcx4fj8Xj/4OBgfzqdTsfj8f5wOBwPBoNEhqfFAAAhhKitJN75eHDOWefcaDwex1mWJd77wWq1Gmw2m8gYkwCIlFKRECLSWscAIgCREEISEZVlKWazmfj0008N0LiK3L26IM+fP+f/8T/+h/feu/F4XCqlMmbW4/F4kWWZrm3pxtba9WazSReLRQYgGY/HGA6HWmt96SoUCLxHmoAuo7bHQquIX7EYQidAfScOXL4sgn2feOdMkJ9sxf0198WDt92OriD1zhvxrgtctf7qWqC0M1w/Tqp5uCqO3pFYQtbH38a27I+GbuCPyMM5B2NMLZJUAkgzz2AwwGAwCAJIIPCBQkRQSrVFxAOBQOAuwszOGFMWRZGv1+v1arWaL5fL2XK5PN9sNqda69dEdKqUOhNCnA+Hw3MhxBJAmiTJ5uOPPy5OTk78119/7Z8/f35XO5UGAreW8KTxy0DPnj0TX375pSAiPRgMIqVU4r0fCSH2vPfTsiyPnHMPjDGPyrJ8VJblI2PMQynlg9FodPT48eOjjz76aPrkyZP9/f39wWAwiKSUMvQ4D/wUCCGYiEQURUoppb33Mk1Tkee5LIpCe++jps6Mcy6y1ioiIq21SJKEhsMhzs7O6LvvvqPvvvsOf/3rX/Hv/t2/w1dffXVnfrSPj4/pH//xH+k//If/QOv1WnjvSSkF55y01krnXMzMMYDEGBPneR4VRaGISCRJIpVSQtyzrl6VVUmK5XKJPM9hjNk6X7gM3U5an2xsCTPf0e/szlxQ7ip34Li4liHS3+b6mK+LUbSvdlzI+PjJaK4xzTDQqcXS8+uvlwCRqAukG5SlgTGm7S0d7LACgUAgEAjcVYwxRZqm6Xw+v5jP5ycXFxevsix7aYx5BeC1Uuq1UupMSnkhhFh471ej0WgDINdam//4H/+j/fTTT/mLL74I4kcg8DMQMkB+fujZs2fiyZMnCoB89OhRzMxxWZYDVMXND6y1hwAOpZSHURQdAZjW4ydJkhxMJpO9Bw8e7D169Gg8nU6HcRzLIH4Efipq7yw9Ho+F1lpJKbW1Vq5WK+mcS7TWI631nhBiIoSYe+/HqOzaoiiKdFEUerlcKinlpizLQkpZnp6emj/84Q/2+fPnwB2xxKrT2f2LFy98nud2MpkUURSR914bYzQRrZxzyyzLFkVRTJbL5SjLsjiKInlwcBAlSaJC79XAbeRtfipu/QnaJfz03Qre1zFzbb1b6tNcn4WvzBv4adlWgLgqiH5pUVZZXFXzlmWJ+XwOYyoBRGsNrS8fSZi5tcaSUobMkEAgEAgEArcF9t43L8/MrQV4nuerzWZzcX5+frJYLE6Wy+WJtfYcwMX/z9697Mh1XXcDX2tfzqWuXd1dTYmSZVtxEoSMkQEFAx5ZGjrzziMkwPcSbL6GH0Gcehgg0igjxYNABJIB4cSMRPalqk6d+9577fUNuqrdbEuUZEtkN7l+QKGr6lQLpwh11Tnnv9da1tolIi4RcZ2m6ZqIqhhjPR6PWyJyABAA4MZ10RDiJpEA5IeFh4eH6u7du3o4HBoiSrbzPoho6Jzb8d7vEdF+kiR71tr98Xh8YIzZAYBpCGGQZdloMpkMZ7PZcDweD0ajUSrBh/g+bebBbBlmVm3b4mw2Q611SkQDa+0UEYfe+2HXdZn3Po0xau+9AgDtvVdEpJIkUUSEs9kMnXPw2Wefwb179whuxvVVBgB49OhR/MUvfhG01uC9R2ZujTGJ1roKIZRd15V935fW2tIYM5jP5zkRUYzxVe+/EEK89uQQ6Hq6Wgnyx4oQvAhCtMaLwcZt2wIRAQDAYJCDMRqc8xdhlbX2ojUWIkovfSGEEEK8cswMRBS996HrOh9jDAAQlFLUdd2yLMvT1Wr1dLVaPauq6lmSJKfGmJW1dqW1XmutawBorLVNmqYtEbnHjx8HAIgffPDBTbhmIsSNJQHID+dy+GG11qnWOu26bhRjHAPAJIQwCyHMQwjzPM/n4/F4/t577701Go12rLXjTWCSpmmazGazNMsyWQInflBKKUjTVM9msxQRJ5uKpZFSyjvnhnVdD46PjxPvfeKcQ2ZWMUaDiAYAtFLKWGs1Iqq6rgEA4LPPPoOjoyM4Ojq69gkBIvLR0VHM8xzatgVrLWituxijRcTaWlvFGEsiqowxlbV2YozplVIkqzWEEEK8ybbhBSJCjHwlDOHnZoRobQAAoe97WCwW0LYdJEkCIQRQSsFwOISDgwPY29u7GJYuhBBCCPEqMTN770NRFO1isaj7vm+ZubXWdkS0aNv2zDn3jJlPjDHPlFJnxpiVUqrUWtdJknQxxq5pGue9d+Px2ANAPDw8vPbXSoS46SQA+YEcHR3h22+/rQDAbOYmZHVdDxBxHELYCSHMAGAPAG5Za+eDweBgOp3O9/b23trZ2ZkOBoMhMys4v6issyzT1lolKx/FD2nTDksPh8M0TVMdQsgAgJRSsa7rzFqbVFVlnHNmUx2hich0Xae11kopZTbPqSzLoK5r6Puef/WrXzEA3Igv9aOjo8jM/PDhQ37//fcjEemiKKy1tlFK1SGEWmtdaa1rY0yjtXaIKAGIEEKIN9q2Fdb2/tb5c+ePt0HG9nXOeSiKNZRlBQAA3ntQSsFkMgGtNaRpCsaYi9+VIEQIIYQQLxkzM8cYmYhC3/ddWZbVycnJqizLdYyxTJKkAoAFES2cc6fMfGqMOU2S5CzP83WapjUzdyEEn6apS5IkAED47W9/KwPPhXhJJAD5gdy5cwefPHliEDEBgIyZB8w87vt+13u/CwD7aZrOsyx7azAYHOzt7e3v7+/v7e7u7k2n0/FgMMgAAJgZr7YTEOKHgohgjFFaawUAZtPTmwEAtNaGiMxsNtMAYJRSuu97G0JIvfeJtdZqrRNjzLY1FmRZBm3b8o9//ON4dHSkbkIVCABs3zMxc/zkk09c13V9CKHtuq6x1lZEtG2B1Vhre0SUfp1CCCHeeFeDj8uBxeVwRGsNzAwxxot2WDFGcM6BUgqICIbDIaRpCgAAw+EQ8jwHa62EIEIIIYR4aZiZiYi8977rum69XldFUSwXi8VJURRL59wqTdOV1nqplFoCwNIYs7TWLobD4WowGNTj8bhVSvnFYkHj8Zju3btHiBgBAI6Ojl7xOxTizSAByA8Dl8ul8t6bNE1TpdTAez8OIezEGHc3ba9upWl6azKZ3Lp9+/Z8f39/NpvNpoPBYGCtNbjpEyChh3jJEOBPengjAECSJHY8HufMzFmWqTRN9enpaVJVVdr3fUJEJk1T65zTxhi1OVDgPM+pbdtw584dukkhCMB5EPLxxx/Huq4pSRKPiD0idkqpVinVGGMapZRTShG/IcN1L6/wFUIIIb7ON31fbGd7IOKmbdYfDw+ICIqiAMTzNll7e3uwv78v7bCEEEII8VLFGNl778uyrNbr9bosy2VVVWcAcGytPQOAFSKuAGCplFoBwNoYs962ziaibn9/v1+v1wQA8d69exFuxoxUIV4rEoB8//Dw8FDVdW2stdYYk4UQhkQ0iTHuENG+UurAGPNWnue3JpPJrYODg735fD6ZTCaDJEkSrbXM+hDXjtbaDAaDTGttrLUGAEzbtrbve9t1nQUAZGYVQgA+L10iZg5t2/pNb8sbGYIsl0s2xlAIIWitnda6Q8QGERsAaJm5I6JARKSUioiIm4szkl4KIYR4422qSS/uA/xpKyyl1EXFyPa5qqrAew/OOUBEyPMcjDEXgYkEIUIIIYT4gfAWEXnnXFOWZXF2dnZWFMVp3/cniPgsy7KzNE2XzLxSSq2YuTTGlMzcAECzXC77uq79hx9+6AEg3rlzR9pdCfGKSADy/cGjoyO8c+cOPn361ACARcTMOTeKMU5ijDve+z1jzH6apnNr7cH+/v58f39/bzab7YxGo8FgMEiVUghy4VRcQ+qc1VobRETvPVZVpYhIIaKKMdKmL2YEgOi99/EDTWcAACAASURBVEopr7X2q9XKv//++z7PcwCAGxWCfPnll/z+++9Ha23o+94DQM/MHTO33vumqqp2sVi0IYRuMBjoLMu0MUZt/paFEEKIN9q2EmQbXFzddnV2SIwRmBn6vocQAgCct9QcDAYAcN4OK8syMMZICCKEEEKI7935yI9IIYS+7/u2qqpivV6frlark7Isj2OMJ0mSPEvTdIGIqxhjEWNcK6UqAGiIqAeAfrFY+J///OcEADIzVIhXTCoNvh94eHio/uEf/kHHGI1zLu26buC9n3jvd733+865eQjhYDKZvLW3t/fWu++++/bt27f3Dw4OZjs7O4PBYJBsWl8hXj07FOIa2P6/qZRSzIxKKdRamyRJtLVWERETEXRdBwAQlVJkjCFEDIgYdnZ2wunpKf7t3/4t7O7uwk9/+lP45JNPrv1BwP/7f/8Py7LUSikTY7QAkIQQ0hhjGmMcOOeGTdOMuq6zzKzTNFWX5qjcaF3XQV3XsF6voes68N5/5evkI0sIIcSLvOh7YhuCXL5t54Nsf8YYwXt/EYhYa8EYA1I0LYQQQojvGzOHEEJXVdWqKIqT5XL5tCiKp2VZPu37/pnW+lmapsfW2rM0TZd5nhdKqXIwGDRpmranp6fOGOP/93//N/7P//xP/Oijj679dQ8hXndSAfKXw8PDQ3X37l09m820c84CQJrned73/YiIpkS0i4h7Wut5nufz3d3d+bvvvrs3m812xuPxMM9zY4y58RdLxZvDGKMGg0FijFFZlkGapuC99yEE6rqOYoyBiPoQQo+ILTN3zrlub28Pmqbhg4MDvn//Ph8dHSHcgP6XSZLE0WhERVH4GKNTSnXOuXa1WtVFUZRPnz5dHxwc5ERkR6ORSdPUWGtf9W4LIYQQ19bl+SBXZo+BUuq5Qenr9Rqcc9D3PcQYIcsysNY+F6xcnikihBBCCPEtMDNv+10BIjIzAxH5vu+b9Xp9dnp6+myxWDxt23bhvV8opRZKqTOt9WmWZes0TaskSZq+77s0TXvnnMuyjACA7t+/H6XyQ4jrQQKQvxzOZjM1mUz048ePE611mud53rbtuOu6KTPvJkmym6bpPMuyg4ODg/ne3t7ubDabTKfTwWAwSJRSUvUhbhSlFFprtdZaISIjYmyaxgFAQEQiIh9jbL33HQC0aZp2ANA550BrzW3b8meffcZHR0d8dHR0rQ8IHj16xLu7u7yzs0PW2tB1nQOA3nvfOeearusaRKy11u3u7m7vnBuyTAkXQgghXuhq6HF1m1LqogokhAB1XYNSCtI0hcFgACEESNMUmBm01mCMgTRNL6pDhBBCCCFeJMbIIYTonAtEFJiZEDESUe2cW63X62dFUXyxWCy+BIAFIq601ktr7coYs0zTtBoMBm2e5/10OnVZlvlnz54FAIj/9E//JMPOhbhG5OzgL4OHh4d4+/ZtvV6vbZIkiTEmr6pqFEKYENEOIs7SNN3f3d2d7+3t3bp169b+pvJjkGVZYoyR2n1x41xqhwVJktjBYJDt7e2NjTExTdNYlqVr27bpuq6z1jYA0LZt22VZxkop6vs+tm0b79y5E+F85s21PjBYLBa8u7sbNzNNnPe+11q3IYS27/t2Mw+kJyKPiATX/P0IIYQQr9p2LsjXrRm4PCidiICIoO97WK/XYK29CESYGZIkgdFoBLu7u4CIEoAIIYQQ4hsRUez73hdF0XRd14UQeq21Y+YyhLCoqur/mqb5ou/7p8aYZZIkhda6AIByOBwWw+GwjTG66XTq27alZ8+e0ePHjyX8EOIakrODv9BsNlNVVenbt2+bpmkyIhqEEMYhhJ0QwkwptZem6Xx/f//gvffee2tvb29vMBiM8jxPpO2VeB1orXWWZenu7i5mWYaDwQCUUs4518QYuxhjTUQtALTMHPq+91VVERHRcrmk614Fcv/+ff7Nb37DMUYiomCtdV3X9YjYaa07ROyUUr0xxm1mnlzb9yKEEEJcF1fDj8vD0re2Acd2ODoRQVVV4Jy7eF0IAYbDIRwcHIC1FqQFpRBCCCG+jRBCbJrGHR8fl8vlsqyqqkqSpDHGLJVSi67r/s8598xae2ytXSVJsk6SpMyyrB4MBrX33uV5Hp48ecKPHz+Ojx494vv37zNI+CHEtSMByF/g6OgIz87OlNbatG2bMvOg7/sJM8+cc7shhH2l1F6McWatnY1Go+loNBrleZ5tWgdJ2ytx411qh5UqpVgpFZ1zfYyxT5IkIGJvjHEhhC6EEJg5JEkSBoNBIKIwm82udRUIIsLHH38c67qm4XAYzs7OPAD0iNgBQGetbTdhiNNae621hCBCCCHEt3D5UPhq+LHdfjUY8d6D9x5ijBBCuKgM0VrDYDC4CEuSJAFjjFSDCCGEEOICMxMRhRBCqOu6KcuyXK1Wp4vFYlUUxcpaWyZJsjDGLJj5GBFPrbVnWuvSWlsBQDOdTtvVatUDQPjtb38b79+/zx988AEAAB8dHb3aNyiE+EpyRvAXuHPnDv77v/+7mk6nxjmXEtEAESdEtOu93/Pe7yqldkIIE2YeWmuzJEmstVb+3cVr41I7LJWmaQIAg52dnR2llM+yLDrneu99771vAMAhYo+IfVmW/uDgwP/hD3+IzByvcx746NEj3rTrouFw6MuydETktNad1rrXWnfW2t5a65VS8VXvrxBCCHHTbI8DrgYhV0OSbUusEMJFCNL3PZRlCWdnZxfbp9MpDAYDCUCEEEIIcYGIqOu6vmmauqqqoiiKVVmWJ03TnDVNs0zTdBVCWFhrV4i4yLJsmaZpYa2tjTHtdDrt9vb23OPHj/221ZWEHkJcf3JG8OfD5XKpptOpds7ZEELqvR8i4k4IYY+I9jcByNQ5N3LOZUSkmfn6XuUV4i+ktdZpmqbT6XSapikMh0NVVVW3Wq26tm1rAGgRsYkxtojojo+P3Y9+9CN6+PChAgB61fv/NRgAcD6fx5OTE3LOBWb2xph+0yO0tdZ2aZp2xhinlIpSASKEEEL8ea4GIds2WZcrQbTWoJQCIgKtNSAidF0Hx8fH0Pc9OOdAaw1JkkCapq/y7QghhBDiGiGi0LZtc3Z2drZcLs9Wq9Vp13XHMcZFmqaLzZDzxWbeRwkAFRHVWuuOiFyM0Z+dndHh4aHM+RDiBpEA5M+DH3/8sXry5IlJ09QWRZEBwCCEMAaAKSLOrLW7SZLs5nm+s7OzMxoOh5k5X4Imcz/Ea0sphQBg0zRVABABIDRNM4sxls65gplLpVSFiI1SymVZ1hMRvf/++5GZGRGvZfXE/fv3+eHDhzwajeJyubwIQTazP1pjTA0AtXOuqaqqMcbkMUaVJIlSSilEvLF/99sLUde5QkcIIcTr5avaYQE83xJrG4xsh6UTETRNA0op0FrDcDgERATn3MXrlFIXc0K01i/vDQkhhBDiZeJ4PsQzElGIMdKm60R0zlVN0yzW6/Xxer0+Kcvy1Ht/YoxZIOLSWrvUWhda6zLG2OR53vZ938UY/Wg08kmS0L1796TttRA3jAQg3x0eHR0hAOjpdGrOzs5SY0y+qf4YhxB2jDG7aZruTSaT3d3d3dmtW7cms9ksT5LEaK3lKqJ4nanNBQYNABRCGDHz1Dm365xbI+IaEUtr7UU7rCRJyDkXASCeZyDX70ACEfno6IjffvvtGEIgIvJaa6eU6tI0beB8VUhZVdX6+Pi4CCEk4/EYJpNJlqapMcbc2AAEQMIPIYQQL9fVAenb57Y/t3M+tuEHM0OMEbz30DQNICJkWQbOOcjzHJj5oiJkPB7DeDyWAEQIIYR4TTEzhBCobdu+aZo2hNDFGJ3W2oUQ1mVZnpVl+ayqqpO6rs+MMWdJkiyNMYUxpsjzfA0ADQD0bdv6d9991z158oQ+/fTTCADxgw8+uJYLN4UQX08CkO+ImeGTTz5RJycnum3bZDAYpE3T5H3fj4hoTERTpdROnuc7b7311s5PfvKT6Xw+H06n02w4HEoAIt4YMUZFRMY5N3DOjZ1zU2aepmm6YuaKmTsAaJMk8TFG+uyzz8K9e/eu7YHE0dERHx0d8WQyIe89IaI3xvTM3CJiVdf1Osa4LIpieHBwYG7duoXGGLW5verd/1581QUpIYQQ4odwdfj59rktrTXEeH7YsH3dNhjp+x5OT0+hKIqL11lrYTgcwttvvw3WWkjTVAJ+IYQQ4jXEzBxC8HVd18+ePVtVVbUOIVTW2oaZC+/9om3bUyJaGmOWSZIstdaFMaZExEopVQ8Ggw4Awmg0Cv/5n/9Js9lsO+/j2l6zEEJ8vdfjqtxL9ODBA7xz545yztk8z9OmaXKl1DBN01GaphOl1DTLsp2Dg4PpW2+9NX7rrbcGs9ksHwwG1lqrNi2ChHjtbQajG2ttnqbpOM/zKRFNEHEcY1xrrZsQQhNCcLPZzJ+dnWk4nwNyXa+w8+eff853797lt99+OzjnPDP3iNgSUU1EZVEU69VqVSDiIMuyfH9/f0BE1/X9fCcSfAghhHjZLs8D+arnroYk24qQEALUdX2xnYggTdOLipAsy8BaC8YYMMZINYgQQghx83GMMTIzee990zRVVVWr1Wp1WhTFWd/3hbV225Vi4b1fMXNhrS2steskSSprbW2tbZm5S9PUTadTOj4+jl9++WX8l3/5F4bre61CCPENJAD5ju7cuYNPnjzRe3t7tu/7LIQwiDEOkyQZWWunw+FwZzqd7szn8+nBwcFod3c3H4/HibVWzqzEGwURldbaZFmWTyaTMTNP+76f9H0/ZuYRANRJkmTW2o6Z+/F43D98+PBaB4QPHz7ku3fvxhACDYdD37atQ8ROa11VVVU2TVP2fV8Oh8NJ0zRdCCEw841eIXK5z/rl+0IIIcTL8lXVIFe3KaUgxnjx2DkHMUaIMQIRXTweDAaQJAkopWA4HEKe54CIF+GJEEIIIW4eZuYYIznnuq7r6qqqivV6fVaW5XFRFMdd1y2NMSulVJEkyQoA1kmSlEqpGgAqY0y7u7vbeu/drVu33M9+9rPw4MEDPjo6kuBDiNeABCDf0b/+67+qv/qrvzLr9TpFxJyIRgAwSZJkuru7u/Pee+/N9vb2dmez2c54PB7meW6l7ZV4EymlVJZlZnd3d5DneRyPx21VVdPFYjEpy3IcQqidc1WSJF3btl0IQc/n8+v+t8IAEOfzOZ2engZjjDPGtDHG2lpbaa0rpVS9CUWcUuq1HY4mQYgQQoiX6Wobxhe1yFJKPRdqEBEgIhARrFYrCCFA3/cwn89BKQWvS6tKIYQQ4k21aXvV13W9XiwWZ0VRnJZleRJCOLHWnhhjzgBglSRJYYwpELFi5kYp1WqtWwBwRORnsxn97Gc/IwCIm/BDCPEakKP9bw8BAG/fvq2ttTaEkIUQtnM/JgAwzbJsurOzM5nP56PpdDpI0zS11mqUBsPiDbRp96YHgwEaY3Kl1JCIRtbaISIOY4yDGGMeY0xDCHY4HKosy6773wrfuXOHR6NRdM4RM/sQQq+1brTWtTGmBoBGa91prR0ixtctAJE5IEIIIV6Vqy2xLg9Gv/rzq76viAiaprkIRKy1kCTJxZD07e9prcEYcxGkCCGEEOJ64HORiGI8HwZGiBiZ2XddVzVNc7parZ4WRXHSNM1pjPHUGHOKiMskSVZa6zUilojYpGnalWXZA4CrqipUVUW//OUvGQD4dTuPF+JNJwHIt4NHR0cIAAoATAghQcRBjHEUQpgw85SZd7TWkyzLRqPRaDAajTJjjH3VOy7Eq4KIqP+IiChLkiQHgCEADGKMA2bOY4xpmqbGOadXq5WC87Dx2h5sPHr0iO/cucMxRjLG+DRN+77vW611AwANIrabAMRrra/zTBMhhBDiRnpRKHG5CuRyUBJjvGiNtQ1AtrNAnHMXc0C2A9IHgwFYa2U+iBBCCHGNMHMMIVDf985774io11p7Zu6cc0Vd18dFUXyxXq9PvPdnxpiFMWaRZdnKWrvedG6om6bptdbub/7mb9znn39Oh4eHr93iRSHEH0kA8s3w8PBQffHFF+r27dsaABIiyohoREQ73vvdzW3mnJt673Nmln9XIS5hZmRm5b1PiCjz3g8QMUfEjJnTEEISY9R5nuPR0RFe91LT+XweT05OorU2eO/dZlBag4gNIjZKqR4RPQC8NgdRX7eaVgghhHjVLrfC2t4/XxT6vG11ByJCCAFWqxV478Fae/EdNxgMYGdn56I9lgQgQgghxPURY4zOOVcURbler6u2bUtjTK21Lpl52TTNCRE9RcQFM69ijEWSJAURVcaYBgDa8XjcTadT/3//93/h4cOH8f79+6/NebsQ4qvJhfoXw6OjI3z77bdVXdfGe2+SJEnbth1sWl/tIOJelmX7eZ7vJUmyo5QawPm/q9TLC/FHiIiKmS0RZTHGnJkHMcZ8E4gkxhidpun27+baVoEcHR3xxx9/zE+fPo0///nPw8nJiVNKdYjYAkDLzC0i9kopj4gRrun7+Lak9YcQQojr7up31dXZIFdbZgEAhBCgrmvouu7iNcwM4/EYiAjSNAUAAO/9cy2yjDEX94UQQgjxw9gMNWciiswcASACAHvv+6Zp2uVyuTg7O1uu1+szY0xhrV0i4pKIzpxzJ5vgY72Z9VEjYuec64nIpWnqnzx5Qo8ePYrwGi1aFEJ8PQlAXmDb9ipJEr1arcxwOEzats1ijAPv/dgYMzXGzIbD4Ww6nc6m0+kkTdNcKSUBiBBXxBg1EVkiSmOMGSJmm1k6aZqmhoh0WZbqzp07yMx8jS8s8OHhIf/mN7+JaZqStdZvKj56Zu4RsUdEp5QKmwBECCGEEC/JNvzYBhpX54JsxRih6zpgZogxXrTIIiIwxsBgMAAigiRJIMZ4MS8kz3NIkkQGpwshhBA/oBgje++p73tHRD6EELTWwXvfNU1TF0VxulgsTpfL5bFSapFl2QIRVwCw1FovlFJrpVS9HXKutXZEFACA+r6nR48ebYecS/ghxBtAjty/Hn7++ed49+5d1TSNGQ6HSYwxd84NQwgj59zYWjsZjUbTH/3oR7P5fD7b29ub7O7u5lmWmc0AaCEEnLfAijGqGKMhoiTGmG6Gn6fee6u1NkSkkiS5EX83Dx48gF/96lf8X//1X7y7u0tEFIjIhRAcETmllNdaB601yWoSIYQQ4uXZhh9XAw+AFw9P384MCSFAWZbw9OlTODs7u3g+yzKYTCZwcHAASikJQIQQQogfEBFR13X92dlZVdd10/d9Y4zpmLnu+76q63pBRAut9ZlSagUAS6VUYYwpELEIIdQxxtYY0yGia9s2AADN5/P46aefxqOjI1msKMQbRI7cX2A2m6nJZKKdcwYAkhjjABGHMcax936MiOMsy8b7+/uT27dvj2ez2SjLMpskicZrvHxdiJdtcxFCKaWs1jrTWudKqRwRU2ZOQgiGiNRwOMT5fH7t/3a2bbCGw2FUSlHf98F7H5jZI6JnZk9E3jkXnHNBa01KKdx61fsvhBBCvM4uhyBXn99SSkGM8bnXbqtB2raFEAIAwMVzg8EAeucgyzLQWoPWGpRSoJSSdlhCCCHE94DPVypEZo7Oub5pmmaxWKyWy2VRVdVaa10rpUpmXjvnihDCSmu9QsRCa10opUqtdamUqtI0bZm5t9Y6IgqTyYROTk74ww8/jB999JEsUhTiDSMByNfYtL/CNE110zQJAGRKqSEzT0II0xjjhIgmSqlxnuej8Xg8nE6nmTq/yvmqd1+I6wa11jrLsmw6nQ4RcRxCWDNzrpRKYozWGKOMMei9hwcPHlzbGSAbfHh4GB88eIC/+MUvyDkXkiTxMUYPAM4516/X6/7s7Kzz3vej0cgPh0NtjNHGGPmAEEIIIX5gV4eiX3V5WLpSCgDgog2W9x6cc0BEQEQQY4TeOVBaw3A4vAg9siwDa61UgwghhBDfA2YmIvLe+75t26qu6/VqtTpdLBbL1Wq13AQdK6VUaa1dA0CptV4rpcokSUpmbqbTaVNVVYeIrq5r//7774fHjx/Hf/zHf7zx8zmFEH8+OVp/MVWWpU6SxHrvM0Qceu/HIYSJ937snBs653IiShBRb1d4v+qdFuK6UUphkiR2Z2dnoLWm8Xjs2rZd13WddV2XxBg1M+svv/xS/ehHP7r2g9ABABCRmTl+9tlneHp6SnVdEwAEIgqr1coBQNs0TbW3t1ft7+9nBwcH2Xg8RmOMetX7LoQQQrwprlZ4bNtgbUOPy4fuWuuL7VtKKSAiYGZomgZOTk7AOwd938P+/j6MRiMJQIQQQojvQYwxdF3XVFW1KopitVqtls65UwBYWmsXxpglAKyUUuskSSpErJm5MsY0WusmTdMOAFySJJ6IwnK5jPfu3aN79+7JrA8h3nBytP41Pv/8c/zlL3+JAKD7vrcxxpSZh0Q0ijGOQwijEMLAOZcRkYkxykVNIb4GIqK11gyHw4G1FofDYb9er0cxxiyEYNu2NQCgrLWY5zneuXPnWocfl/C9e/diWZb09OnT4JwLMUYqisK1bdudnZ3VZVnWRDQcDocmz3P5zBVCCCFesm34sb0PcF7tsX18uVpEa33xWGt90SYLAKDvezg7OwPnHIQQIEmSi3ZYl+eObGeKyLooIYQQ4k/wZkECb1peXdy8923btsXZ2dnJarU6LYrizDl3ppRaDofDpVJqYa1dMnPJzI21tmHmJsbYd13XI6InIsrznE5OTvif//mfo8zkFEIASADyte7evYtffPGFstbqyWRimDmJMeYAMGDmQYwx995nIYSEiDQzyxmOEF8DEVFrrZVSyhjDWuvcOZcZYxIAsDFGo5TSWZapJElwPp/j17WsuE42VSB8cnISm6aJcN6vNLRtG5qmcTHGDhH76XTqvPcUY5SDLyGEEOIV+KpjiquD0rdVIVe3aWMuBqRvZ4MgIgxHI0BEcM5dPKeNhizLILEJWGt/yLckhBBC3Dib2VpERME552OMAQCCUir0fV82TXNaluXT9Xp9UpblmVJqgYgra+1q0/6qSJKkjDF2aZp2Ozs73Zdffunfe+89f+/ePQIA3nx/y7m3EOKCBCAvMBqN0Dmn+r43zJwgYua9z0MI2/DDhhBMCEHHGDHGiFrrV73bQlxHuLmQgACgN2GIiTHaGKNhZm2MUVprfPLkCQLATZgDssXL5ZIBIG5v3vtIRBRjDM654L0nIpKyWyGEEOKauFz1cfnxV23btsFCRCAi8N5DXddwfHwMdV1BmqQQOYLWGvI8h93dXdiZ7oAx5tov5hBCCCFeMg4hhKZpmqIoqr7va2ZujDEdERVN05zWdX3ctu1ZCGGRJMkKEUulVGmMKbXWlda6zbLM5XnunHP+7bffDr/97W/pgw8+iK/6zQkhricJQL7GF198gTs7O+icU0SkEdFYaxMiSkMIKRHZEIL13mvnnHLOYQgBEJEvrRiTMx4hvsKmYgqZWW3mfygiUlprNMZgkiR4//59ODo6etW7+o0Qkf/t3/6Nz87OuO/7bRXIcz/hfBWKhB9CCCHENbatPt2GHZdtj++3bbF618NyuYT1ugCA85ZaSZLAeDwGpdRFBci2FRYzX9yXUEQIIcQbYNPhCratrgAAOMYYnXNdWZbl8fHxYr1eL0IIa2NMiYirGONZ0zRnIYQVIhYAsGbmGgCaEEKrlOryPO8RMcQYQ5Ik4fHjx/Ho6EjOt4UQX0sCkBdo2xa994qZtbXWIKJ1ziUhhCSEYPu+12VZ6tPTU3z69ClorXk0GuFgMIAkSeTkRoivwcwYY1TMfHELIeByuVTvvPMO3rt371Xv4nfy6aefAgAwETEislIqMnNUSkWlVERE6T0qhBBCXFOXq0AuD0y/GJy+ed3lY/tIBE1TQ9wMViciSJMEQggwHAwhscnF/JBtcJKmKSRJIpUhQggh3gQcY6QQQnDOBWYOcL440LdtW1VVtSyK4mS5XJ72fb+y1hZa6xUiLpl5xczrGGNFRFWapq3WulNKubqu/a1bt3xZlnE8HtPjx4/j4eFhBOm2IIR4AQlAXqDve0zTFBFRMbMmIrtp2ZPEGE3btnq5XOLvf/97JCJomobfeecdODg4QK01GCP/vEJ8nc2J/0UAopRCpdTF1YCHDx8iM+NNCA7u3LnD//Ef/3ERgFwSt4PdNoPeXvWuCiGEEOKKy0PSt7aPmRng0nBz3gxPjxzP+5gTAcUIkSI48NC2LSxXS2BmKMsSAM5baKVpCtPpFCaTCSCinCcIIYR4rcUYOYTgy7Js6rpuvPcdIvYA0Pd9XxZFsazr+rSu67O+71dpmq4Qca2UKrTWa0SskyRprLUNEfWTycTFGMNoNCIAIADge/fuxXv37km3BSHEN5Ij729ARKi1Vt57HWM0MUa7CUJM13W66zrlnIOzszNeLBZMRJjnOQyHw1e960JcW5daxKHWGhERY4xqNBqBtRYfPXqEh4eHr3gvvzutNYcQtiW+l1tgCSGEEOIa+6oQZPv8pQcASgEwg0YNFAm01oCoIGIERADvPSwWC6jrGrTWwHwegIzHY3DOQZIkkCTJS3xnQgghxMsXY+Su63xRFOvj4+NFWZYlEdVa6zrGWPZ9v2rbdoWIS2PMmpnXWusySZISEWtmbvM8b2OMfZIkbrlchvl8Hk9OTvjDDz9kkDbTQojvQAKQr7FcLvGdd97B7XDzTRWIIaLtTTvnVAgB27aFruvAWgvvvvsu9H0PMco1TyFehJlxO/tjMxwd+r7HxWKB7777Ln7yySf44Ycfvurd/FYePnwI77zzDiultre4GXq+bXy6Lcm9sQdoUsEihBDidXe1LdW2DdalJ57bfh5wMCAyaK0uviudc+C9B+DzShGlNFAIkFgLg8EAmBm2LXO11qCUehlvTwghhPjexQ3vPW0ppWKMsa/rel2W5fGm1dUqhLDWWpfMXALAmojWAFAkCz7e5AAAIABJREFUSVIBQJ2maWOt3Q5E7wHA/f3f/7178uQJffbZZ/H+/fu8+V6WE1MhxHciAcg3ICI0xmwv0urNwGYdY9QhBOWcwxgjAgBUVQVd1wERyYVCIV5gE37gdhh6CEEZY1AphQcHB696976zu3fv8mq1AgCAEMJ2eCrzeQ8vBjgflv5Kd/J7Ip9tQggh3iRfGYIgXFx6QUA4zy8QODIwwsVMEIDz4egKI7RdB+uyhPTsDIgIQggwmUwgTVMJQIQQQtxYMUbu+57quu7atu2cc84Y0wNA23Xdqq7r46ZpjruuWxBREWNca61LrXUZY6zSNK2UUo1zrlNKdUmS9G3b+q7rwv7+fvjd734XDg8P40cffcRHR0ev+u0KIW4oCUC+hRgjnofYSsUYNRGpzQBnBAC8dDH3Ve+qEDfC5fBjM+cDN+3mcLlc4q1bt171Lv7FNlVg23ZY8uEghBBC3FB/cozPz7fMQjifDwIaAK600trODAFmqKsKiAi6tgXvPVhrwVr7kt6FEEII8f0joti2rT87O6vPzs7Kuq4ra21tjCkRcdG27anW+nQwGCyZuQCAQilVMnOllKqTJGlijD0z+7IsAwCEp0+fxjRNY1VV8fDwML4uiwmFEK+OBCAv0Pc9fkXI8dzK9W31B4CsjBbiz3Q+Df3SAPQnT55s219dWmN5c2wO0KQnqRBCCPGaunzcj5eGpAMA8HZg+maA+vb1fd+DDwEQAOymHVaMEdI0BWYGpRRorcFaC8YYqQwRQghxbcQYIxHFTZeryMyEiNE519d13RZFsVoul8uiKNbW2tJaW1hrl8y8AIBFnucFM68BoMyyrHLONczcDAaDrus6n2UZ/eEPf4gAEBeLBUu7KyHE90kCkBdwziEiotYaAJ5ftQ7nocj2eQk/hPgLaK3BmPOPo/39fUjTFD777DO8d+8ebCpEbuQfmMwCEkIIId4MF9UgiBfBBcJ5GAKbcwUiAu89VEqBsRZskkDTtmA2s0SSJIE8z2EymQAAyLB0IYQQ1wYRxa7rfFVVnXPOxRh7rbXz3jdN01Tr9XpVFMVitVqtkiQprLXrJEmWSZKsh8NhoZSqjDF1kiRVjLGdzWbtarXqlsulPzw8DIj43MmztLsSQnyfJAD5yyAAPLfiSwjx3SilbmS4IYQQQghxeUbIxeKo81lgF9uuhiPBe6jKEmKMsF1oFYlgMBzC7mwGWmvQWksAIoQQ4togIqqqqnv69GlVlmXVtm2VpmmFiKX3vizLckVES2ttoZRaA0CptV4jYk1Etda68d53zNxaa5333hFRAAC6qQsehRA3hwQgL5AkybZ//1fanOzglcdCiG+AiH/SHsoYw2maXjx379697fDwl7173xtpXSGEEEK83i4HHQDwXOiBiH9SDbrd1jsHYROUxBghxghd3wMiQp7nAAAQQrhojaWUAmMMGGMuQhMhhBDie8YxRiaiGEKIzBwBICJirOu6q6qqXK1WxXK5LKqqKtI0LbTWawBYO+cKRFwZY0qtdcnMdYyxYubWOdeladolSeJCCH69Xvu+78NyuYxffvmlhB9CiB+cBCDfglKK6fwE5eKi7eUe/9L+Sog/DyJyjBGYmb33AACwu7vL8/mcAQAePHjwSvfvz8XMqJTCEMLNTW+EEEII8a09N/j8SuXH9qdS6rx1LgB478F7fxF+EBHEGMEYA1mWARFBXdfAzGCMgSRJYDgcQp7nEoAIIYT4QTAzhBBi3/e+aRofQnDM7JVSvuu6Zn1uWRTFqizLpbV2aYwpjDFrACiVUmulVKW1rpVSjda6ISIXQnBFUfjRaBSIKFhr6enTp/HLL7+ko6MjBpnzIYT4gUkA8i1dDj6UUrwJQ7bbbvQqdSFelc0FgucOdk5OTqAoCnjy5Mmr2q3vFZ5/OMgHhBBCCPEau9zmCuB8Dtg28LjaBgvgfP7Zdpva3DhGaJsGjp89g+ViAUqpiyHpo9EI3n77bWmNJYQQ4gfDzOycC6vVqnv27FlV13UVQqiNMS0RVV3Xrdu2LZi5yLJsZa1dWmvXxpiSmStmrrTWDQC0Sqkuz/M+hBC89wEACADiF198EWezWfzyyy9Zwg8hxMsiAcgLpGnK3vuLD+Nt1QcAsFKKtdacZRlba2E6ncJsNoPhcAjGGAlEhPgOlFJsjOGmaWA2m13dfO0PiD7//HN85513AAAuhrl77xHPS8Tkw0AIIYR4zV2dA3K1AuRPKsY3oQcgng9K3/y+cw5CCBe/H2OELMvAOQdZlv1J+LFtjbWdGyKEEEJ8Rxxj5BgjhRBCXddtWZblYrFYrVarwnu/1lqXiLiOMa6dc2tEXBtj1tbalVKqSpKkYuYGAFpEbBHRIaIDAJemKR0fH8fZbBZ//etf84MHD+Bf/uVfJPgQQrxUEoB8C0op3tyi1pqVUhEA2FrLWmve2dnh+XwOt2/fhp2dHciyTHr/C/ENLrWU403bBx4MBs8dBN2/f5+Pjo5e0R5+N1mWYYwRQwi4aYF10febmSUIEUIIId4AL1oEta34uJgRsqkQgc1w9E3rEdi0BwUiAiIC5xwwMwyHQ7DWgPcOYuSL8CPPc8jz/GLIuhBCCPFtMTMTEXnvXdM0bVVV1ercYrlcnnVdt9JaLzftrQprbam1LrMsK5VSpTGmGQ6HTdd1fYyxR0Q3GAw8EYVf//rXAc5niEjYIYR4pSQA+Ra2La+01oyIUSkVlVIxyzKeTCbw/vvv449//GN877338Pbt2zAajWQFlhDfDm/byr3qHflL9X2PSikEeC7wUCjlYEIIIYTYuFwh8lUD0lGp54aoa61BKQUhBFgul9D3HSRJctFiazAYwnw+vwhDJAARQgjxXTAzbwaT14vFYlkUxWq1Wi1DCAtr7SkiLhBxoZRaGWOKzYyPSinVEFGjlOq99/35fyaE+XweTk5O4nw+3w5Qv/Hn+kKIm08CkK8xm80YAEBrzUTExhgyxgSt9fZGaZrG2WwWf/rTn/Jf//Vfw7vvvovD4RClAkSIF9tWf2zDD6UUb1aecAiBb1pv67t372JRFEBEaIzBrwLnc0AkDBFCCCHeQJdDDYBLbbEQLw4QcNsSaxOSbOeEAACEEKAsS6jrGgDOq0OMMTAej0FrBUmSgFLqYhHW5ZZbSqmLbVpradUrhBBvCD4Xt5h5G0hsz8cjEVHXdXVVVauTk5OT5XK56LpuEWNcWWtPkyRZGGPOmLkwxhR5ntdKqTaE0C0Wi56I/Gg0Cm3b8nw+jycnJ/zo0SO+f/8+S/ghhLguJAB5gaZp2BjDWZbFTeVHMMZ4pVRARErTlIbDIe/t7cFbb72FBwcHqLWWMwohvoVN+BG11hERo9aa8zzn+XzOy+WSP/zww5tysIQA5y2wiAi89yrGqGKMCgBw+3Pb8kIIIYQQb6arxwEXc0KuHCNcXUi1nQXSdR2ctw2liwDkvDXWCLIsByJ6rgp9G7IYYyDLMsiyDAD+OK9MCCHE642ZYwiB+r533ntHREEpFZRSpJQiRCRmdk3TVOdjPxbPiqJYhBBWaZoWWZadGWOWWuulMWY9GAzKJEmaNE1755ybTCb+ww8/pK8KOm5KK2shxJtBjn5fIE1TNsbELMtIKeVjjM4557TWvbXWWWuD1po2F3BvysVaIa6D7aqTGGPcBiCRiPiLL74AAOCHDx/C4eHhK97Nb8bM8Jvf/Ab/+7//G2OMatMGSwGAZmYNAIqZlcwAEUIIIcRVl4elXx2kfnn75fkeiH+s6giBYL1eAzPDcrl87r9HRMDMkOc57OzswHw+B0SUAEQIId4QRBS7ruuLoliv1+uy67pGa91rrZ3WutNa9wDQOeeq9XpdhBDOAGCNiGtErJi5YOYKEUsiaoiodc65qqpCURQE5+f0r/hdCiHEN5Oj369x+/Zt3lSARK01MXMwxvRJknTe+15r7Ywx3hhDWuu4mRPyqndbiOuKNwM9mS5BRNJa0yYIYSJi5xwnSQKHh4fXvmSWmfHBgwcIAJgkCcYYlfdeG2M0ABhEtFmWWWut3gQj8iEhhBBCiD9xOfQAeD4M2YYafwxAEM7XkgDEGKGua/DeX2yPMV7ciAjG4zEQEWRZBlcrUrdBitrMHhFCCHEz8B/7W23vXrSa3t53zvVd19XL5XJ5cnKyKIqiMMa0xphGa11rrVutdUNEVdd1pXNujYiVUqrRWtfM3CBiG2Ns8zzvy7K8GHA+n8/jp59+yrD9QhJCiGtMApAXGAwG7JyLSZIE55xXSvWI2CVJ0hpjemOM31aBXPcLtUK8SpuTcOr7nvq+79u27Zumcc65EGMkpVRkZq6qCv7u7/6Of/KTn9yYv6c7d+7gaDTC3/3ud2q9XisAUKPRyGRZlmRZlh8cHGQ7OztpmqZGWuQJIYQQ4qqvqwK5Ojdku/08rADYZibOOXDOAcAfww9mhhACEBGEQKC1gTzPIYQAbdsCwPmMEWPOn0+SRCpDhBDiBiGi6L2nrusCEVE8b0dAABCNMQQA5Jxrq6oqV6vVycnJyelqtVoqperNrUTEWmtdA0CNiI33vt6EHa1Sqh8Oh53W2uV57gEgJEkSxuMx3bt3LwJA/Oijj27MebsQ4s0mR7lf45NPPoEPPviAR6MRAUCw1jpE7IwxbQihsdZ2SZL0SZL4bQusTQgiFziFuIKZue97Wq/X3Xq9ruu6rrqua9q2dTHGYIwhpVSczWbx97//Pfz+97+HGzIDBOfzOZ6cnCgAUIiolFJ6MpnYg4ODbH9/f7S7uzva29sbjEYja4xR3/hfFEIIIcQb53IIcvX5y9svV3Bsc5HLv7sdcr6dB4KIECNBXddwfHwC63UJ1hogIkjTFIbDIczncxiPxxKACCHEDRJCoLIs3WKx6Nq27Z1zzhjjtNZ+07GkDyE0fd+XbdsuYowLAFhrrSulVG2MqbTWNSI2McaGmdvhcNgqpbr2/7P3LruRXMn9f8S55KUuLJIS1aI0Y8mC4QW1lOGNF5IAw4ABb+VHGK/8DF16Aq+tR1BvvPDKK2k7xsDwQlz84P9gBtOj7uatqvKeeS7xX1RlMStZxe6W1GqyFR+gWHk5efJkVmbyZHxPRJRlEwRBY601ZVnaLMvcaDTycRy73//+9/TJJ59wGHiGYe4V3MvdwdHRETnnPAB4RGwFkNI5V6wEkFIpVWutjZTSCSH8624zw9xViIiMMTZN0+r8/DxPkiTz3heI2CilrPfea629c45+9atf0ePHj193k59Lm9NjPB7jn/70J0FEQkopm6ZRe3t7wYMHD6Jf//rXo8lkMhyNRnEYhooFEIZhGIZhdtH3BOlPd8WQ9rsftqq/jbUWiACqqoKrqytYRuRc5gcZDAYwmUwgiiJQSq0TqLd1tgIKh8ZiGIa5ExARrUNfVVVl0jQtnz17li0Wi6Isy0IpVUopq5W9KgeAfBXeakFEizAMM611LoQogiDItNblys5VKaUqY0yFiM3R0ZH505/+ZOu6dmEY+idPntB3331HH3/8MU2nUw57xTDMvYMFkFuYTCYURZFDROOcq+M4Lowx+UotL4IgqLTWtdbaCiH4HwDD7ICIyFrrq6pq0jStFotFCQB1FEUNItogCFybBL1pGjo/P7/rOXXwyy+/xE8//VSUZSkmk4kYjUayLEultZZRFKnxeBwcHByE4/E4iqIoEELgHT8mhmEYhmFeM7sEjXa6nw+k3aYrkAghgIjAew9KKSACcM5CURhYGc/AOQfGGAAAmM/ngIhgrV3Xp5SCMAxBaw1a61d92AzDMMxzWD3XnXPONk1j0jQtkiRJZ7NZMpvN0qIoUiFErrXOpJS5UioFgFwIkRFRRkSZ1roIgqCI47gMgqAkogoAaillU9d1E8dx45yzH3zwgc2yzJ2enm4IHo8ePXqt54BhGOaHwgLIDj7++GMCAF9VlTs8PDTOuUpKmWmtoyiKBs65NIqiPIqiSill2AOEYW4HET0RWedc7ZxrAKBGxGa1zFlr/WQy8WVZ0unp6Z0XFE9OTnA8HmMYhuLq6koJIbQQQgNAgIhaSqm01lJrLdjzg2EYhmGYH8I2QaQreHjv12W89ze2bcv2hZTWO6QoCri4uICyLCEIAiAi0FpDGIZweHgIe3t7oJRiLxCGYZjXD1lrbVEUxXw+z+fz+fzy8jIpy3JhrV147+dCiMRam3rvUyJKEDFDxAIAiiAICu99LaWsAaDWWjfWWjMYDEyapu74+NienZ2577//3v/TP/2TW9nE7vx7OcMwzIvAAsgOHj58SF9++aXf29tzzjkDAPVgMMi99xERJcaYLAiCIgiCUkrZGnH9ynW8HenNbwoMAwCISEIIL4RwUkorhGgAoEFEo5QyUkprrfXWWirLsu1k3dnO1nQ6xdPTUxyNRiKOYymEUCvRQxORJiLlvZfeewH8HGAYhmEY5iekFTO6IshttInT2+2892sPEmMMzGYzSNN0LZYEQQDD4RCklKC1hiAIbggg/TBcLJAwDMO8NLR6LtNKzKbVwvU0AKynvffeGFOmaZqen59fXV1dXS4Wi0Vd1wshxDyKoplSao6ICyFEopRKACCXUhbGmKqu6zqKoibPc+u9t2EY2vF47OfzuX/nnXd8mqaUZRk9efKkzW97Z9/HGYZhXhYWQHaAiPD111/T06dPvZTSHh0d1U3TSGNM7pzLgiBIhRCpcy4tyzItiiJVSkVhGAZaayWEkPwiwDAbkBDCSikbKWXtvW+EEA0iNgCwFkAAlgLkdDp9zc29nePjY3TOyTzPNREFRBRqrUMhRLiaV0Qk2lwhDMMwDMMwPxVdEQTgZs6Qls2k6csybW6PNhRWWZZrIcV7D0EQgLUWhsMhKKXWgkk/UXtXIFFKbYTlYhiGYW7He0/ee9c0jbPWWu99m1uWhBAOlgKEb5cRkc3zvMjzpfPHbDa7zPN8gYgJESVKqZmUch6GYaK1ThAxI6JiOByWRVE0qzBX9uLiwv/FX/yFOz8/p3/4h3+gL7/8Eh4+fEgAsCG8MAzDvEmwALIbOj09pePjY39wcOCaprFBENRCiFJrnWutU0RcGGNms9lsjIhR0zR6f39/NBwOB0EQcMB/hrmGENELISwiNlLKWkpZCSFqIYRRSlmllDPG0Pn5+V3vdCEAiF//+tfCGCOdc7ppmkgIEXnvYyllREShc04T0RtjCegaPBiGYRiGuVv0Q1wBXAsh/QTq3TBaba6Q7jcAQFmWMJ/PAQAgz/Ot4bTCMITRaASTyQSEECyAMAzDvATee1/XtU3TtCyKomyaphFCmFXEBAMAVghhV+/QlohMVVVFkiSLPM9nRVHMm6ZJV6HaU6VUgoipUipDxFwplYdhWAkhaq21KcvSAoD713/9V98XOu764EOGYZgfCwsgt/Dw4UN69OiRBwCX5zkGQYBRFFXe+yIMw9R7P8/zfPj48eN4sVjoPM8lAIBSSiulNL8EMMw1rQCilGqEEBUAVFLKWgjRKKUMIvooivz5+fnrbupzOT4+xj/96U/y/fffV9baoGmaGBEHSqkYEWPvfUhEGgDeqBBYLIIwDMMwzP2hK3xs+x/eH6ullALnHCAiGGNgsVhAWZarROrXHift9Gg0gqOjIwjDcO0FwjAMw7wYzjlfVVVzdXWVnp+fJ2ma5u0gwfYbESshRNPm7bDWFmma5nmeZwCQImKBiIX3vnTOFWEYFgBQCiEqa23tnGtWIafd6emph+XARH6pYxjmFwf3Um8BEWk6nRIA+JOTEzubzQAAaiIqgiBIrbWzpmnCsiyDpml0EATR22+/HXvvR4joAUC+3iNgmLvBKgeIk1I2SqlSa10QUaG1LqSUFRGZuq6dEIJOT0/pLjtPffHFF6KuazEcDuWTJ0+CKIoiIhoQ0ZCIRt77ofc+cs4Fzjl530JgWWvBGLM2fOR5DsaY58YXZxiGYRjm7tFNkr4tRFZ/fpXPEIgIqqqCpmnW61rxoxVWrLWglII4jsFaC2EYbuwHAEAIAVJKCIIAtNbr+hmGYd5knHPeOeeapnHOOU9EbWgrj4geEX1d13We5/lisZjNZrPZYrFIhRAlLAcKFohYCiFKRKyklJX3vgKAsmmasq7rkohKpVRlrV0nNldK1d77ZrFYGCmlmUwmVkrp/uM//sO/9957fmXfYhiG+cXBAshzmE6nNJ1O/enpKZycnNimaZq6ritrbQYASVVVUV3XkRAiNsbsEdEBEVkeKc0w1yAiIaJf5f+opJQlEbUdupqIjJTS1XV91xOg48cff4zWWlHXtdJa67quIyIaWGuHRDQAgAERRatk6PI+hcEiIjDGQFmWkCQJzOdzSJIEmqZhAYRhGIZh7in995LufDc0Vn+d9x6ccxvCSTdMlpQS0jSFq6srqKpqw1Ok7TdorSGKItjf3wdEZAGEYZhfBM45l+e5ybKsquvaWGsNIrrVoEArpTTGmKosy2wVzmpWlmW6Ej0KIUQBAMXqfbkEgMo5VxFR5ZyrEbFGxFpr3TjnTFEUNo5jAwCmaRqLiM4Y48qy9Kenp342m9FXX33Fic0ZhvnFwgLI86HpdEq07M37f/u3fzN7e3vVaDTKsyxLvPeBcy4KgmAYBMGh1roSQjh2K2SYa1YjBb2U0mityyAICmttIaUstdYVETXee/fkyZM7Pyrl+++/x+FwKOSy1xqscn8Mvfcj7/0IAAbe+9g5F3jv75UHSCuAJEkCz549g/l8DkVRQF3X65AYLO4yDMMwzP2k6+nxvJBYbSjfVvRop6WU63nnHOR5Dt77dfirrpeI9x7iOIbJZAJKKVBKrb1EGIZh3mSapnFZllV//vOf0yRJyqqqylV+j0YIUSulKkQsnHN5lmUJACziOM4QsVRKFYhYSClLAChXYbAq733tva+dc7UQwlRVZZqmsVEUWWOMn8/nTinlhsOhn81mdHBw4E9PTwkA4NGjRyx+MAzzi4YFkBekFTT+/d//3e7t7TXOuSoMw8wYE0opY0QcEdGiruu0LMtMCDEIwxCUUlIIwQnRmV8ctMQ757wxpq7runTOFQBQSClzIiqklKVzrgYAo7V2H3300Z3umE2nUwQADMNQWmsVImrnXEREQ6XUeG9vb288Hk/29/dHw+EwVkopIcS9ufeJCJxzUFUVpGkKaZpCXdcboz0ZhmEYhrlfdJOed2nFjTbBebusm/AcYCmGdD1EunkOjTHrQRIAsJFQ3XsPdV0DEcF4PAYp5XpdmzRdaw1KKU6gzjDMfYScc9SGu1qFufKI6PM8L9M0zRaLxfzq6ioriiIXQlRSykopVbUiByLmxpgMANIgCIpVuKtSKVUKISoiquM4rowxzSoXSGOMMdZaK6W0w+HQPX361Idh6K+uruiDDz6gVvT4l3/5l7seXYFhGOZngwWQl4MODg58nud2OBxWRJQHQaCttSEADMqynC0WiysAOKjrOhyNRjQajWKttZZS3hsjKMP8FBCRt9a6uq7rqqryoiiyqqpS730qhMiCIMiklK1bb5PnuYc73jk7OTnBPM9FWZbSWqu896H3fiCEGMdxPBkMBgeDweCto6Oj/f39/VEURVrcozf61ihhjIGqqtaxv1sjBcMwDMMw949d47C6SdK7y7rb9AWP/jrnHBhjNjw/+rlCpJQwm83AOQdZlgERrfOCjEYjGAwG7BnCMMy9g4jIOefKsmyKoqibpjGIaIQQpiiKLEmSNE3TWZZlaVEUKSIWQojWuyMXQhRa61wpVSiliiiKSgBolFJ1EAR1K3g458xkMjHOOfPOO+/YxWLhJpOJOzs7899++62fTqccq5hhGOY5sADyknzxxRf+q6++csPhsAnDsKzrWhtjYu99OpvN5tbay9FoNDk8PAzeffddDIJAKqUkALD1kPlF4b0na61J07RM0zTNsmzeNE1irU0BIFt1/kqtdW2MMWEYusePH99lAQRPT0/x+PhYeO9FXddaShkQUQQAw9FotHd0dHRwdHT09sHBweFwONyL4ziUHOyaYRiGYZg7Tt87pBv2qjvdLdcVS7aF1+omS5/NZpBlGWitwXsPWmsYDAbw4MEDUEpBEAQ7hRqGYZi7yGrgmE3TtDo/P0/zPC+896UQorLWplVVJc65eRAEKSIuiCgXQuRCiFxKmSNiW74UQpRN0zRCCBNFkXHO2TAMbZ7nTgjhyrJ0i8XCn5+fu6OjI39ycuJPTk7o888/v8vvzwzDMHcGFkBeEkSEr7/+2ud5boMgaJxzlRCiWLktLuq6nhVFcWmtjbTWKoqigIgwDMNQay04HBbzJtMNe1VVVVMURZVlWZokyaIoirlzLkHEDAAKrXURRVEVBEHjvbeHh4f+v/7rv+5sB246neLx8TEeHByI77//XgVBoOq6Dp1zcRAEQwAYDQaD8eHh4XgymQzDMIyUUpK9vxiGYRiGuS9s8wDpr+uzTQDphtSy1kKWZUuPUkRw3kMYBFDXNaxCBt/qjdIihAApJWit2TuVYZhXChF57z0555z33nnvCRH9KjQ6IaJfeX9UWZZlV1dXiyzL0qZpCq11QUSpcy51ziVKqVQIkSBippTKvfdtkvNSa122eT2klGYwGNgsy/zR0ZHLssyPRiN/fn7uZ7MZPXnyhL777jv6+uuvPcB1mHaGYRjm+bAA8vLQ6ekpHR8fu+FwaIQQtbW2MsbkTdOkzrl5WZaXRBSFYRhEURQ653Bvb4+Gw2GotUY2iDJvKkTkjTGuLEtbFEWZZVmeJEmSZdm8qqo5Ii6CIEiFEDkiVt77GhGbX/3qV/bBgwfu4cOHNJ1OX/dh3ICI8NGjRzgajUSWZTIMQ1WWZUBEgXMuMsYMAGAopRwMBoM4juMoCILgdbebYRiGYRjmZdgmfLTLu+JIX+To0k2g3obXtNYCEIEnAvIemiAA5xzEcQxCCDCNAehU0w2j1c4HQQBxHMNwOIQgCFgAYRjmlbGKZmDLsqzVExJcAAAgAElEQVTruq6NMVZKaYUQDhEdIjrvvSmKokySJF0sFvPFYpEaY3IpZS6lzKSUGSJmWutMCJFqrXMiKrTWhfe+stZWzrl6MBjURVGYPM8tAPjZbEYA4AEAfve739HDhw+pK3bweFqGYZiXhwWQH8DDhw/p0aNHHgBcWZbWe19LKUtYhvWZI+KwLMvw2bNnsqoq8dZbb7kHDx5Mjo+PcTweCykl99aZNxJrLZVlaa+urvLZbJakaZp47y+89xdSykul1FwIka68pqogCJo8z20URQ7ueP6Pjz76SDx58kTOZjNtrQ0QMXTOxU3TDLz3g6ZpImNM4JyTRMS9UoZhGIZh3hjaZOkAuz1BWvrr10nYYalxoBBA3kPdNHB1dQVFUUA7bqQVTNp9tvNEBKPRCA4ODuDdd9+F8XgMSvGrLMMwr4aVd0d9fn6ezGazJM/zQkpZK6VqKWWNiA0i1tbaMk3T3BiTAEAuhCillOVqwF8ppSyJqACAAgBKAKibpqmDIKgR0Witm6urKxNFkfnjH//oT05O6MmTJ/Sb3/yG2mfudDq90+/JDMMw9wHuNf4AEJGm0ykdHh56pZQ1xjQAUCFiLoRIAGBQ13VgrVVFUQTeezkYDNTR0VFERDwqnHljWYW/MlmWVfP5PE2SZB4EwUwpdRUEwQwAEkTM4zguiKgCAKO1tkVReFi6Et/Fzh0CAJ6dnYnFYqGCIFDOuaCqqtA5F3nvI2NMZIwJnXPaey9YAGEYhmEY5k1im/jRenjs8gbZlS+EAMATgbUWiryAuqpBCAEE114f3vv1p022XlUVAAAMBoN1bpJtnipCCFBKgZSSvUQYhgEAAOccOOfAWnvj2dF9fhERSCmttTYpiqJIkuTq/Px8niRJqpQqhBDVSuSoELEioqJpmsIYk61yeVSIWK9EkBoRKyll7b2vVwNnTdM0xhizzvURRZEFAPfw4UO/asudjIrAMAxzn2EB5AcynU7pN7/5jX/vvffs4eGhQcTKWpsTUeK9D+u61mVZKgAI4zgO6rqOrbUTet6QKYa5xxCRt9bauq7LoiiyPM/nRNQKIFeIuFBKZYhYKqVq773Z29tzf/jDH/zHH398J+8NIoJvvvlGZFkmEFESkXbOBQAQElFkrY0AIGqaJjTG6DfFA6QbdoJhGIZhGAbg+QJHt9wuT5B2nXMOvFt6e3TFD4ClsbIVQtppRAStNQyHQ/DeQ1VVa2+RFiklKKVgOBxCFEUsgDAMA7QSXKuqgqIowBgDzrmN/EXdbyGEEUKcZ1mWLxaLq9lsdjWbzRarBOZF+1FKlYhYImJBRKWUshJC1ADQKKUaa60JgqCRUhrnXPtxo9HIXlxcuMVi4ZqmcQcHB/6LL77wd3QwIMMwzBsBCyA/HJrNZv69997zzjmjlKqVUgUipsYYrZRSRKSFEIMgCIZKqYlSyvI/NeZNBhFJCOGUUlUQBKmUcq6UulJKXUkpZ0qpBSJmQojKe99ore3l5aX79ttvPdzREFhffvllm/xc1nWtAEBLKQMiiowxkXMuWk2Hzjnlvec3bYZhGIZhfhFsS14OAGthortu23RXEFmHyiICIcTaA0RKuZ4uigLOzs4gSZJ18vR2X22ekNFoBEdHRyCEAK31qzx8hmHuAUQEdV3DfD6Hs7MzyPMcrLXr50/rOdZOK6WKMAz/v7Isi6IoFog4D4IgW+X2KIQQORGVSqlCSlkiYgUApXOuRkQjhDBaayuEsHEc2yRJHBE5KaWfzWY+z3P/xz/+0QOAb5Oas52IYRjm1cICyI/g448/puPjY2ettURUa60LRJRKKcBlr14JIWKt9QAR96y1edM0sVgihRAIAGwsZe41tMR77721tnbOlVLKVCm1CIJgprW+1FpfrLxAEkTMiahsmqY5Ozuz//iP/+j+5m/+xj9/T6+Pg4MDHI1Goq5rZa0N6rqOiCgKgiAWQgyEEMPBYBBrrUMhhEDOTMcwDMMwzC+AfpdnZ/6PLUJJd/R1a3zseoEIITbCYRERVFUFzjmQUq7DYAFc5wuJogj29vZAaw1a6w0PkG4Yrm6oLPYSYZg3hzbUVVccdc5Bnucwn8/h/PwckiSBpmk2RI/utJSyCMPw/znnyqZpMkTMwjAspJQFIhZBEBQAUCJiFUVRpZSqnHOVMcZYay0AuMPDQ5dlmb+4uPDD4dDPZjN6//33CQDo9PSUAK5ze7D4wTAM8+phAeRHMJ1O6euvv/Z5nts0TYX3vtJaIwBAHMeSiAIhxAARh865SVmWiyAIQkSEIAgiRFSIyD1u5l6zyvvhjDFNWZZl0zQZEaVCiIXWeq61niHiXCm1IKLMOVchYuO9N3Ec3/nk5wAAo9EIZ7OZVEqpqqoCAAiFENFgMIiFEMMwDIeHh4eDwWAQKqUUCyAMwzAMwzBLWuGhK4YAwIYwcptI0i1rrQVr7YZQ0k2UbowBAIDxeAxhGG54h3TFGaUUhGEIcRyzCMIwbwhtyLy6rqFpGjDGACKCcw7SNIUkSSBJElgsFmCtXd/3fRGEiEpE/L0QopJSVkqpIo7jSkpZaq1LRCyDIKgBoJZSNkKIOoqi5v333zcffvhh+357l3NcMgzD/OJgAeTHQV988YX/6quvnLXWHB4eQtM0BADgnBNKqUAIEVtr4/l8HgFAUFWVm0wmZn9//wARB0op/g2Ye41zztd1XSdJkuZ5Psuy7KIoiivn3ExrPZNSzhFxEcdxUtd1EYZhZa01k8nEnZyc3Hl335OTE3z27BlOJhORZZkCAE1EgVIqmkwmg4ODg/H+/v7+ZDLZOzg4GAwGAyWlZAGEYRiGYRimwzbvkP60935DJOknWO+LJ22ZdroNl5UkCTjnNkSQ1pNECAFRFMH+/j689dZbEMcxCyAM8wbgvYe6rmE2m0GaplCW5fr+r6oKsiwD7z0EQbDh8QFwQ2wtEfGPiFgDQO29r4moMcY0iNggYgMARmttmqaxw+HQGGPs5eWl++///m//xRdfELD4wTAMc6dg4/uPBBFpOp264+NjMMYQEdFgMKA8z0UURQEARM65cD6fB3meq6ZpBBFhGIYaEeXqI3DF6z4ehnkRVmGvCAC8tbapqqpIkmSepullmqbn3vtLIpoFQTBXSi201omUMg+CoPTeN4PBwD5+/NifnJzci07hcDjELMukc061CdCVUtF4PB48ePBg+ODBg9FoNBrGcRyFYagEv0UzDMMwDMNs0L7qdEWNrojR0k9s3t2+b6zs1y2EAOccZFkGVVWtw2i13iOtADIajdYhs6SUNzxEurTtFUKsP/zaxjCvnm4IvG5eoe692vUeM8ZAnuewWCzg4uICiqLYEEBbD7HW62vbc2gVWq+SUv6ZiBpENABgAMA652xRFC6KIuucc3VdOwBwQggfx7H7z//8T//w4UMWPhiGYe4gLID8BEynU5pOp+7TTz+l8/NzX1WVt9aKKIqUECKo61qVZSmapgFEFFJKDIJAO+fAew9hGIZSSiWllK/7WBjmRSAib621zrmmKIo8y7IkTdOLJEnO8jx/ppQ6C4LgIgiCmRBigYhp0zQFADRBEJjHjx+7zz777M57fwAAnJ6e4kcffSS01qqqqoCIQiFE1Ob3GY/Hg4ODg8FwOIy11gG/EDMMwzAMw+ymb3Rsp9ucHtv6Uq2Q0a+nn0y9rauua6iq6oYB1Tm3NpQqpSCKIrDWrpOlbxNCiAiklKC1hjiOIQgCYCd+hnn1OOegaRqoqgqMMeCcA4CbofHaeWstZFkGs9kM5vM5FEUBzrm1h1f7HGmFzJauB9qqvmZ/f//ZYrGwRORW4Z6d1tpHUeRPT0/p5OTEz2YzOjg48L/97W/p4cOH9Pnnn9N0Ov05TxHDMAzzgnDP7aeBptMpTKdTf3JyQvP5HN999926aZrSe58KITQRKSGELMsymM1mEgBknufu8PDQ7+/vTwaDQcwCCHNfWI14qbIsy/I8X2RZdlVV1RkRnQkhzhHxUggx894nWutcSllJKU0Yhvby8tJ/9tlnHu5B7g8AgOPjYzTGiLIsFSJqa23ovY+IKCaikIg0AMhV7nNWPxiGYRiGYV6AbUJIy7Y8If3tttXTTaS+zbukLWuMgTRNQUoJSZJseIp0t21HjwdBAMPhEI6OjmA8HrMAwjA/A+19enV1BXmeQ13XG2JGS1/8TJIE6rpeCyat51dXYO3nJOp6mACAzbKsFEI4772bzWZeKeXfffddms1mBMv3WHry5Ak9efKkHRB7L95tGYZhfqlwz+2ng6bTKRERfvnll+7dd99tBoNBmWWZDsNQOuekEAKrqtLOOZFlmcjznLz3QmutpJRSCKGEEAgAbEhl7hyrkFdERGStbcqyLBaLxTxN08ssyy6cc2fe+zOl1LlS6lJKOZdSJt77ommaOgxD8+GHH7o2Mdx98P4AAHzy5AkeHx8LrbWy1mrnXOici4goWgkhGgA45BXDMAzDMMwP4LZwWH0jZXd5v45dIay6o8XbcFfOOcjzfO0J0m7fDbXTjgYnIojjGCaTCURRBFrrtQBy2z77iZUZ5pdIe78B7A5v19IXOquqgjRN4fz8HBaLBRRFsRGGblv+DuccGGPAWrshpHZphZB+ezrip9daV0+fPvVhGPokSei7776jjz/+mACWEUDaTX7QSWEYhmF+dlgA+YlBRCIi9+jRIyGlbCaTSVGWpYiiSBRFgc45Xde1ICLhvRdBEOjBYKCFEEhEEIZhwOGwmLuIX2KbprFlWeZ5ni/yPL8qiuKiLMtzpdQZIl6EYXiBiFdBEMy11mkQBGWapqabFO6eiB8wnU7xgw8+EHmeK+ecJqLQex8BQOy9j733kbU2ICJBRG/km+02YwTDMAzDMMzPxbZ4/93lrUjSDaG1rd/SD5vTNZJ2jaGtEHL97aFpagAAmM/nIIQAYxoAwBtiTbc9SikIggCiKFrnHGCYXxLOObDWQl3X0DTNOgfHNi+ubV5ebT6PJElgsVhAWZZbxcW+ENL3IGs/3fu8+6zoP2Occ3R0dGQePXpEX3/99Tps86NHj17JeWIYhmFePSyAvAIQkb7++muntV72jAGgqirQWkNd19Jai957LMsSZ7OZkFJCXddmMpmYg4MDDofF3Emcc7YsyypN07woinmWZRdFUZwbY86llGdCiDOt9YUQ4goR50EQJGEY5nVd18YY83d/93fuk08+uS/iB06nUwQAIaWUYRi2+T8i731sjBkIIYbGmNg5F3jvBazu9TeJbclKGYZhGIZhXhfb+iRd42Z32a5tutNdY2i3ru7HewJjLBRFDhcX51CWBURRtPIWoa31CCEgjmPY39+Ht956CwaDAQsgzC8O5xyUZQmXl5drD442B0c/f09XzGjX1XUNeZ5DURQbYiXAtVDZFz/a6f59vyuJei/0VbsdffbZZ+7zzz8nfgdiGIZ5M2AB5BXxxRdf+G+++cYBQJNlGRIROudAa60AYO0BMp/PZdM0VBSFrarKh2EotdZiVa4NhcX/dZnXwdq113sPxpimLMv86upqlmXZZVmWZ4h4jogXURRdSCkvpJRXiDhDxNR7n0dRVI5GoyZNUwv3KOzVdDrFk5MTBAAxm81UXdeaiAIiigAgBoChEGIAADERBQDAgiXDMAzDMMzPwC5xo+uBsctrpG907Sdd7woh7Xy7D2MMzGYzSNN0nU9guR7Ae7f6Xm4vpYTxeAzOORgMBhthtjZB6NtXu23l8FnMXaPrIbXt2uxe403TQFEUcHFxAc+ePYPFYgEAm6JHe413BZB2eetB0jQNAMCGJ1Vf8NzmVdK/v7vld4mmrQByT95bGYZhmBeEBZBXRBsK65tvvgFYChhtbg8VhiF679E5B957qKrKAoDVWrssy0QQBE4I4bXWgRAiEELw78S8Frz3zntvrbW2qqokz/N5nufneZ6fl2V5NhgMzoMguFBKXWqtr6SUcyFESkQ5IlZKqeby8tJ99tln/r50IlvPj6dPn8r9/X2ltQ6stVFZlrEQYqC1Ho1Go/FgMJjs7++P4ziOV/coD+tjGIZhGIb5mdll5LxtfStGtMnP22WtcbUfQgdgOZq9KMq1YLHMbbAMkbU0qF4LJm2ukcFgAEmSABGB1nqLWAOAuPwGoPW3EAKUUhCGISilOOk6cydo82u0Cca7OTRa8aJ7X5VlCWmaQpIk609bti94bPMCaYXG9n7ph7zaRV8E7S7f9b1NCGUYhmHeHLgn9QppRZCvvvoK33vvPby4uAAhhMjzHKSUnoicc841TWPKsjRFUZgkSbyUsiKiZjAYTMIwHLMAwrwmyHtv67ouq6rKsyy7LIrisq7rc+fcGSI+W3mAXGmtZ0KIWSt+KKXKpmmaDz/80H744YceEe9LLxJPTk7w6dOnsq5r5ZzTABB572Nr7TAMw9FgMNh76623Dvb39w8PDg729/b2hkEQKOTheQzDMAzDMD87L9oF2zZifFsOj13bXQsc14LHUrRop69ZeU9DnudweXkJZVmCUmpjv214LUQE8gQE18ZYrTVEUQSTyR6MRiMWQJg7QXtNLxYLqKoKjDE3wlZ1Q7215YuiAOfchtDgvV+Xdc7dECO35fZ4Efr38fPmX7Z+hmEY5n7CPalXzCofiC/L0r799ttgrQXvvZNSNnVdN0TUBEFQSynrqqqqs7Ozumma0hjTICIqpSKlVPy6j4P55eG9h5XnR75YLC6SJDkriuIcAM611mdKqWdKqfMgCGZRFC2IKFsJH9Xbb7/dHB8fGwC4V+LHdDrF09NTeXx8LMMwVGEYhlmWxUQ09N4PhRDjvb29yfHx8eHR0dHb4/H4MI7jQRiGWkrJPWeGYRiGYZg7Rldw6CdC38Zt4bOkFEB0LYjsCq/Tjl4vyxLOz8/XIbC69bc5RIhoKYC0oggRRFEEe3tjQAQIwxCiKPrpTgjD/ECapoEkSeDp06eQJAlUVbXVgwMANkJY1XW9zovTCh1dwQPgZgLz7rIut4W4uy33D8MwDPPLhgWQn4F//ud/9l988QX8/d//PR0cHNDh4aFzzhkicojojTFOCGGdc/VsNmsQsZZSNmEYIiKStbZeJVmWSikppdRSSiWEkDzqnPmxEBH5ZZwr5723zjmPiA4RTV3XWVEUl1mWPSuK4llZlhdCiAut9QURncdxfKG1XgwGg5SIqsVi0Tx48KA5Pj62AODukfjRIhaLhYyiSE8mk3A+nw+996OmacbW2j1r7R4i7g0Gg/F4PB7t7e0NlFKhEELwvcgwDMMwDHM36SU43uoB0q7vbtPPMYIo4Dqq6+bo9G1dQWPMOgTXZo4SAKKVAOLpWgiB5XQcR+CcgziOQSkFxpiNNm1jezif1li8aVxujdVSSgiCALTW7GVyz7HWgjEGmqZZh6fq5765bRrg5v3RJ01TmM1mMJvNIEkSqOt6az6PrvfGMlScA0TcCAPX3ee2/XfZJXJ0xU2GYRiGuQ3u5fw80KNHj/zHH39Mf/3Xf01lWfooijwAQFmWGAQBVFVFq1wLLkkSJ6X0URQJIjJZlmXeew0AYRAE8Wg0GkRRNNBas9GV+dEQEVlrbVmWdVmWtbW2RsRGCFEZY5KyLC+KonhW1/WZ9/5SKXWllLqSUs601gutdWqMKRCxaZrGPnv2zP7qV79ycJ1E/V4wnU7x+++/x/fee08qpXRd1xEiDpxzY2PMnjFmz1o7ds6NAGAQBEGotdZSSn6OMvePH/miSMDhAhiGeXk2DFevsR0/NfxMvD90jbK7jLxdo2o3nM912U3BozX63hRLcG2EbnMKtGJI6/0BAOBdO73KI0IEiMt65/M5AABkWbbzmJYhua6TPnf3D9AJs9UzNF+H2ZpwmK03gG54qrqu16JZS+tx8SKhpbZ5SiEi5HkOSZJAnudQ1/VWAaS9Z7qeHt029Pe7Tdho5/v3VLd9twmBL5InhGEYhvllwb2cnw+aTqcwnU79p59+Cu+88w6dnZ1hFEVisVjgqrPgnHPeGOPzPDdPnz41s9ksJaIDa+1ASjkaj8f777777ltSSqW15sTLzI+GiKhpGpskSTGbzdKyLDMAyJVSGQAsiOjSOXcBAJdBEMyklHMAWCilFgCQB0FQWmvrwWBggyBwn3zyiQcAwnuS9LxLGIaiLEsJAMF4PI4AYFTX9cQ5t++cmxhjxsaYgbU2sNZKamMgMMwdpm9w/MkuWh5txzDMS4I7pn/62m+h/+zaMJL9iOda33i3sQvuLtw1+kbVbflButxWblsekb4BuS+QLA20y/JCChDi2uArYCmGNE0Ds9kMiqLYKk4sxQ5a19N6kSzb4Tfas/Q42TQ0x3EM4/EYADjM1ptA0zSwWCzgz3/+M6RpClVVbQgQXc+MvkCwTRBpt+tet62HSdM0QEQgpdwQAvsCxy5vkts8r7aFwGqFvb7HxzbvEX7eMgzDMNtgAeTnZS2CPHz4kM7OziwA1GEYYhAEZIxxzjnvvXdVVTWrPCCFc25hrR0HQbBnra0Gg4EPw9AjYoOIGgDQe7/2BiEisfpGIQRKKYVSSkgpERFZMPkF4b1vw1t5770nIkLEVpygVYg1W5ZlmWXZIk3TeZ7nCyJKgiBYKKXmRDQTQlxJKWdElCilEkRMtdYZAJRCiGYwGNjLy0v3+9//3n/yySf+PoofACD+8i//UlRVpRAxqKpqAABjpdRESnkYRdHheDw+mEwme2EYxivPD+5hM3eL5RDQtSEOEQHb5QDX0225DrddzP0bGpeV8w3AMMyaFw5BsuX50+fFn04bFb9QeYRNI/VyelfbacvU9jrbZ2JbW7tsvX1/n2ykuxPsMpb2xY2u4bWd7o5s79bXL/ci+27/dVPHu8R7B1VVQdM069H01Pl/vjIBr8WOpbdJu4x6hmKAvuE4jmPw3sNoNIIwDG/NrdBus+ucvej9v200/4vS3aYbvktKCVLKl67vZVjlRlx/nHPrdS9qcH+R8/ZD6mqvtSRJYLFYwGKxgCRJoCiKraJHX+zoeob06+57jSw9l5bnol2/y5tk2z3Qv6daj6ht56JbplvnrnPGwgfDMAxzGyyA/PzQdDqlhw8f4meffWb+7//+jx4/fuxns5kjIiOEMN77qqqqwlpbeO8zIpo55/a01vtSyiJJkkZrXTVNM0bE0HuvvPfSey+JSBCR9N4LIsIwDGUcx3o0GgVBECh2bf5l4b33TdO4LMuapmnMKt+MX33cyuvI1HWd53k+z/N8VpblzHs/d85dSSkXSqm5lHKulFqEYZgppfK6rkvnXDEYDCqllPnDH/5gv/32W//w4cN76fkBy/dIEYahtNZqa21ERIPVfXcYRdHR4eHhO/v7+++8/fbbh6PRaCil1ByCjrlzIIKAlVFkJXSIzvTaA6QngjzPM4R60wgIQH6rQXD9Irtt4x/IC99qW/d1Hx9Jrwq8dfbHwjG47xa4/vNivMrfb6MZSyvvc9u2a/W25Zttv71iIlqXuA5dtT3pLt0igGzuEZdGaEQARLg2USP4lcCyrrXz7OU75u5xmyDSnd4lbtwWtme78RbWF8K1cbrNEULrMEbr7W54GrV1boob/Q/AzRwK7Qj+q6srQEQoimJdb9cw3T+Ofh3983bb6P7nCSDPE4xaY3gQBOvwXXEcv3IBpE3k3QoLdV2v23Rbe2+jHy7teXVtK9e9DrMsg9lsBlmWbW1jP0F5vx3bPEK2zW/zEukv794juwTBbji4Lv0y284FwzAMw7wsbA1/TSAiEZH/q7/6K/s///M/BADOOWeMMSaO4xoRK2NMBQBl0zQ5AGRKqdwYUyVJUlprEynl2HsfE1ForQ2893r1Uc45BQBiNBoFb731ViyEQCGEUEq92t4hc6dwzvmyLM3V1VWRJElVVVUthPBSSiOltIhohBCVcy6v63ouhJgHQTBHxHkYhpdSygUiLoIgWDjnsrquCyFEiYjNYrFonj59auI4dt9++62fTqc0nU7v47s8TqdT/OCDD8R8Plfe+4CIIufc0Dm3J4Q43Nvbe/v9999/55133nlnf3//7eFwGEdRpIUQ3ANn7gRdwxoRgVi9IJP3gK0I4v3SHLcWQ7AdCg0rSWNZ140XS+r8vd5ju/SG4LGqY5sA8kMfED9UAOkbNpnn82OM4HdJAPm5Hs67jnj7XfTy/JjjeBkB5Kf47frh9jancWP5UizYVnrbko6RcMt+r+vseYC8gN7XlTdWA+d7Akj/76bjRiugLB+jy2cqIa1FkJXZGYCuhRFqH73ddrBHyL3hNg+Jbpl+2J+b4sdKNAOEbf+qNkflL5Ovt6JI90pZl0G6sY/l/HbhpRU/jDEwn8+hrmvQWt84xm3TfaGlfy5uE4u2nbNd+9v2v781iA8GA5hMJiCEAKUUhGF4o+xPibUWiqKA8/NzuLi4WOdkuc37oC9W9K+JfniobSJD19OoX65fvmkaqKoKjDEghACt9Q2BYpuA8iIiTtuONqdNO73tWLZdB9vmX2YZwzAMw/xYWAB5jbQiyOnpKX366af+/Pzcee+d995qrc1gMLDOOSOlrL33FRFV3vs6TdOiLMsEEUfOuYH3PnbOhd770DkXEJFeJU1XdV2HUsrh3t5erbWOpJSaiHDVOVnbu9o2tct6nTXstPnW5bQjJ0K7z9vYte22fb/MdneVvqfEFnfeXb0/6pdZdTjb5WsvjLquTVVVVZqmaZIkRZZllRDCSikbrXWDiDUiVlLKzHufAECitV5IKRda65nWeoGIqZQyQ8Q8iqLKWtsEQWAfP35sAcD99re/pel0enN4zj1hOp3i8fGxLIpCSSm1MSYkotgYMySiMQBMpJT7w+FwfzKZTPb390daayWXQ83u5bXHvFnc8OogAlyJHXI1LQAAvV+uW39Wz9Utozc3n7c9oyKtTIUrYx4C7hY/VqNYbzS4V/Nzj/F5hkG6bfaHvUjflxGGL2co2HFM+NwSP+p62JgAACAASURBVHE7ns+LtmPXyP8f++u9jHR2yyW+s8zLtOPHlHlh7ZBewCVj13679/StIshNx4/1fndegxuVb1nfXbdlTUcL2XqNbhm13hdAqCOAdEVVos7zDhEIEQgQUCB4AAAhgLCdXo2ExqVHyFo4aY2F3VHx9+TZ80tlm6fDNq+PXeLINe311q18c+La0L307RQCgehm+EmCzX23l1ErfnTb2p92zq29BaSUW8WNjX3d4tGya5uuJ0B3urvutv1sO+dtfou9vb21cPMqKYoC0jSFxWIBs9kMkiS5IURsEzNuW9dlmxCxzdNiW5m2bu89OOfWwkT/vCDiWlhr6+xOt+3cRl+s6R9b/7fd5unTX/b8e4RhGIZhfjpYAHnNrAzVBAB+Zch333zzjUuSxO7t7dk0TS0RNWVZ1kRUeu/LNE0zIpp774fe+wERxc65iIgi732IiAEAaO99AADRYDAYZlk2UkpFABAAABKR8N7jSpXA1bINQaQrlHS/d61rl3fr6JbtiS7dcwBEhNvWbRNkdpXpsi0m7/P4qYWUXQJGb7RMv8yGuLESyTbKruapc+208361TZuE3FdV1ZRlWZVlmWRZVuR5XiJio5SqpZQ1AFRCiDIMw0xKmQkhMq11qrVOgiBYSCkzIsoBoHjw4EGZJImJ49icnZ3509NTv/L4uM89Vzw5OcGnT58K55wiokAIERpjYiIaGmPG3vsxIo7DMBzFcTyM4zhCzqXD3BV6xsZWCJEAIJwH9A6EJxDer4SQpUAiCAC8B4EI4Gk9Uhw7Rpcbxr71Pq5HNi/HNl8b8zaMiau2rA2E1C7f7jVyG9fld2xxiwCyXcx58X2+3FY/LzeE8xslXvDfWqtt7TBev0BDXn6fz+FFarlpOPmBAkjXOt/b9kV++zspgODN5TfOF+6cubHdlg7arXW0gsOGbRevy3SNrNhp7Dbxo61n+TTaFEG6e9x5vFvrXpUB2Hg+tcrXenbtyXH9HLxxzKtnHyECoQASq2nvgYRYfjyBw+X2AgFc57j8SryhTpgs6jaKBZF7wy6RYRcbRmW8+f/qer5rRF59r68Z3PhfvVnvTQN8P+cCIq4TW3fbvU2s6K5v6+ou7xq+vfc3jOrd/e/yFugb0bcZ0tt5rTUsFou190O7fb/cy7Br+7IsIU1TSJIE8jxfhwvrCwLddvent9XfXXabANKfvm2/AJvhrrrb0Mp7ozvdP9ZtYse289/f//Ou/9vqYBiGYZhXDQsgdwhEpOl0Sp9++qnVWhMAkLWWiMgQUU1ExcpAPXfOxYgYSykj732slAqJKCSiUAjRTgda69AYEy8Wi8gYEwZBoGmZI0QSUZszRAghkJbJ05GIxKqT1IoS608rmLTLe+vF9aGsxY51mU59G2JKt2y7bjUiZfMVc4sI0/3ul215nrDRr++noite9KB2fbdcK2isXgwIOiJHt0xLK3QAgAeAdU4PAHCI6IQQ1lrbVFVVW2szrXUZRVElpWy9PipELBGxFELkiFhKKQulVBGGYa61zq21lbW2DsOwvry8bD755BP7zTff+M8++8x//vnn9138gOl0ih999JGoqkrleR5UVRUS0cB7P7TWjqy146ZpxnVdD40xgfeehQ/m7tB9vqy8OpYeHwTCOxDOg/QEwloQzoHwbimCeAJBtPIKWb0w0zJsFkDHtreeXxpmuoa/9a6xDf2yml5t1q5f2/CwXbFccC2ubDEe3yo87BgdfYsAsmvpbcL687bubvqzPgRvHUy8a+ULHCfeOnurkeJ5osu1QXcz78IubhjNt5XZusft+91W/62npGfX33lWEeFGr2GbJnBLHZsVPr+uXb8D9gv2quwLAdt2ujZ83da0zjOC2ht/ObNRsv+bt/cLbZS7nt4QM7BT93KrjXa0IgFu+dXbZTeMcNgvt1nztufUWmxtn3Grfa/P0vqZ2HqALIUOkAI84kr4QCApwQsCJwikEOCRwK0MkR6W4odYGb89ARAs94fd/dB1W5g3j21G5m0CQbdMd70Hv/H8J2r/D2/PudBnm8F+W5luW1tjd9dj5Da6hvbnle+fg+5+uyilwBgDV1dXUBTF2tvhVQkg1tp1iClEhCiKtpbtelXcVveu37gvCvXFkf6yvvDRLdMt238udoWoXdv1Ba7+9C4Bi2EYhmHuIiyA3DGm06mfTqcAAPC3f/u3YK0FrbUjIhOGYQ0AJSKGq0/gvQ+JKELEQAgReu/D9rtdZowJ0zQNqqrSSillrdUAIIlIrr4FIgpcjmpvBRDsT7ffcC127CoLbbmuiLISWNbCSk94WIsetMWrpDuahTpeIbTDc2SXqNGf74162dpj+xEduY3eb08N6Yog1Fm/Fj1WIsda6GjnYSmSECJ6IvKr9Q4RHQA4KaUVQhgAsETUOOdqIiq01q3o0UgpS0SsiagUQpRCiBIAqiAIKkSsvPe1tbYaDofNYrEwjx8/th999NFa/Fi1+V6LHwAAJycn+Pvf/15JKdt7KUbEYRAEIynlHgDsjcfj8WAwGCqlQkSU3euRYV4bHWNlG9Jq6eVBS7HDOZDWApql+CGdA+EsoGs9Qq5FEEEACKu8Iavq19f4yhiIiKuwV6tddx/1awPgpiGxb06llVUGVwrJjQcibH/edl65V+3YUvYHCCAvxY120ZapF6lmt2HpheuA7SEjdj+VXl4A6S7a1b7dBnPcMtU1mq+2f4Gm7DLst9tviiXb97uxTfdYblFWXlTAwM61v2vb59WxWeHudtwqfvRmbv3Fr9WMjd9wwwC3cx+4NqxuLMX1I2nDENvtEK49KDZs+WtlpNss6J6I7m+8fixtbNcVQnot7wg/fWFtXWTjQFfPOYLr3xXaa627rPfMw2WoKxICSMrltJRAUoCTAlBIQCmBpASLACBWcfiFALESQkgIaCUW6j5Xe+KHb4+D+yFvNF2jctew3Ddat+u3GeJf9n9Lu4/+9C6De79Md7ttgsltfefbhJ5+u1raHBRt+K7bknH3672tHbu2JyJwzoG1dp1fo9v22wSHbe26rS27BJDb5rvbtuv6ERF2/U637bsvfPTFDxY+GIZhmPsCCyB3kFYEybKMTk9P6YMPPrBSSjkcDmsppUJEHcexstbqqqoCRAyCIAgAICCiQCkVOOdCRAyFENo5F6RpqgBAEZEiIg0AsvtBRNEKGCshRMBKwFglel7P08prZFV27TnSEUi624JzTnSFkK5I0hEdul4fa+GjXd9x1cXOCKIN8WOb6NEt772/0TPr1rXr9/gxHbpOp5DaUTRCCGrnsRPmaiVqtEKHx03vD98RUNr5tecHADgicohohRAWEQ0iGillAwCNlLIKgqBeeX/USqnKe18jYtV+vPeNc64Jw7AhImOtNXme27feesuVZem+++47Oj09pTfB8wNg+Zv/7ne/E//7v/+r4jgOiCgGgKH3fqy13ovjeBLH8eTg4GDvrbfeGsVxHEopJXfwmddN+1LaJjMH70EQAVi3FDicA2wMgDEgrAU0BtBaAGPWHiDo3DJMFq0e2ADLOhCvhZCOWLE0ti0Nc23IjdZA146C7gofrUiyFk5gZbhv5zbtpxseIVuPuV1/y4v2NkHl9hP5IoVgfew/tpqfir6xeofp98UqeoHVNw0k7f9av6Oam+1pf67bBJBt+7tNALltf322Gpm2qBy31vG8ZrTVPuc6flGeJ0B1y6znegLIiwlBm0LIbfvo3gnL67C3rl8Pdn+d1lDWbSRuih/9irGzHrvnBNajcdYLrmWRrVVd77ZnDF0vvRZlb4oiK8MfAFDb14SVQZoAQAgARPBCAEi59ABRS8EDlQIv5fKjJIAQgHJZ1qMALwQIgeD9MlzRMozWdTsIr/fpYfO3pfWzmXkT6Ysb2wzS3bItfYGkW6b/fNo234osu8SObc+4fvnb9tVft2t+17O0W957v/bIaNc9T2x5EWFi1/qusV9KuXNQQ/8YbmvT8wSF7nz39+mX2bZu23XR3c9tQtFtbeuvYxiGYZj7AAsgd5TpdOqJCB89egRHR0f+/Pzca63ROeeklNZ7LyeTiXTO6SAItBBCSSm1c06vRBBNRAEiKiGERkQF14KHcs6txQ8iElLKtQdHV9yAlWDRFzradc45IYRAKWU7De26VszQWmObb4R63h7QETtWYsR6vj0XfRFDCLHhCdIub6f769rpZc7qzWXPyxVCLzjaf5uAgps5O0ApRZ3l6+mVMELee1iJHCSE8KvYua2nR1cMWXuA+OWJ9Xjt/eGEEJaIbOsJgqucHwBghBCNlLIJw7A2xhgpZU1Ejfe+EUKYIAjswcHB/8/eu/RIclzn3885EZGXunb1bdgUCQmCYNgt7wh4ZUNaGP4v7O3oCxjw12D31/DeG883eFejvQkvDBGGIAs0IJCUKHnEmenuqsyIOO8iIrOya6qvM+Tczm9Qk9l5jcysazz5nKddLpdhNBr5P/3pT+EnP/lJ/Ld/+zf59NNPJZ+Ld0L8AED/9V//ZS4uLorz8/OR937Stu1cRHaqqlosFovFgwcP9vb39xez2Wy2s7NTlWWp75nKa6X/UY11ByCJACH0YgeaBmgayKqBtC1i0yQxJAsgwQeYGNEXNhCkbBCshY+uU63vruxEAEn167tuxE4ISW3LEslAQJFBOzfH+51nbvNee90yL3TOXrf8Hd/FrsweweUO4ps2e1MHyLXrXjl+u86HG0WAK5pwlcABxEEH9PXr9Id9i878rce59RA3Ooeu3PIV+90igFzHbbt4Xnln0BXOhX5/g/+Hozet0z8f8uv1qufg9qnUCxKy4cJYX+oX200b66+XGXbi4YXxzQOiLJy8uG26tN8NKQ2Q+MLxJGfbppg7CClHJ+rKuuRVFh5iPmLp3jMN95kfsAYwBrC2H7K1ENuNG8TsGOmG0oknXYZI3kcnhBCSCAJan+m3/guZciXbOs+Hwsa2ju77CiHDecMSTlcJLtvaOPz7KpFkW7s3hYLN32bXCSvbRKHN7V3V5pu4i6hy231cJ/5sExQ2r8NVwtBV533bc2DznNzlOXWbY1QURVGUNxXtzHuDyR3lUURwenoaP/30Uzx+/DhMp1Oaz+f83//936Ysy2Y2m5nnz5/bsixNFjosAOu9d8450zSNzUPD6VuladvWxBg5QzHGXvSg1LNOmwDop+f2deIGbyyH4fLGGAy3B6yFjG5fQBIouvFN1WG4DPKvPmsttq07FDquWL//+zoBZCiqbNvmtuWugpk7MUS6v7vxTugIIUBEJC8rIYR+ORERa23sRJJuurW2F0BijNFaG6y1IYQQrLXeWuuJyItI65xricgXRdESUVuWpWfm1hjTXlxc+PPz8/DRRx/5o6Oj8Nlnn8Vf/epX8fPPP5dPPvlETk5OpCvN9raThUV+8uQJW2udMaZqmmbsvZ/FGHdEZGGt3R2NRruHh4eLw8PD+Ww2mzjnjLVWHSDKa6V//nWdfDGmElghAM0KWDWQ5RJYrYDVCmG5AjcryKpBbFtE72FEICFCILBIThKJ607k4TOcaeDikCx7UK5RT5eXJlxeeShAUHcHONZ3b/f3Xt/wmupFjevu6Lzh7xtXuGYx6sSfWy7/XXJJrxjc2n7vd6UbBJDt2+162AcdTnJFR9OWP24j9mzb0NVCzM1T+87rqxa+Y5OuFReu6vi6YvwmtgkJ17ajf81df66vuja37Bq8JFhtEx+2Cze0sa9OLL28TQzEj+6dY5sWslUfGQhiMnScXFru8vPhUqdfX/8KW5aR/r2v24uwSaJHJ1wYBtgkBwgbwCUBhKyFOAd2FuRcGrcGYizEWsAlp8haEGEIMSIn0UNAiJ0IEqU/8b1Ic5/XlfJWcBfhfLPzfFMY2BzepnP/2s/ejU75qwSTbdO3uQlus97mvrcd49AJcV8299s5+bcJMduWv6q9Q246L9umbV6321y/2+zjuufOtmUURVEU5W1DP8XeQmTtnKDPPvuMnz17ZqbTKdd1zRcXF6ZpGuO9NyEEE2M01lq21nKM0XjvuXNtdKWpunFgLTwwJ03De0/deDe/Gw8hdGIGb5tPRNQts0UcwXA8hEDWJj1uc3zz+O+y7JDhfjth5jquE1Su2u5VdAJICAHGmF4M8d4j76MXRIbDgWASN6d3GGOEiIIxJmbnSCzLMnSh6J0rxFobjDG+KIrgvQ9VVYXRaOR3d3cDgIAcpp4fXd7IO8VQ/CiKwpydnY1jjDur1Wo/hHAYQniwWq1+8ODBgx8cHR19fHx8/MOjo6Oj2Wy287rb/n3gvce3336LL7/8El988QW+/fbbvq7yZnjltjvGlO8HAlIHYS59xd6DmgZ8fg66uAAvl5CLC+D8ArRcgpYr0GoFtA04uz9YBFZSFogTwIYAJwIjEb0sTIRtEnF/lzQ2bsIePg+GP6Q3exM3BIXbCiC34VadzHfY4LptL/92+CreUK8SQLbNv1Ubrjm8a7pT+pW2nZ6b23BLMWlr58uWdtzF3HHnE3Q1d3nXu/Z5ecsN3UkE2XhOXNr/jU6g25+EywLE5c6z27RtqJpeel4MO/sGI1sFjy1/D4WY7YczfMIOimINxvuhbJbGyu3lFHbu2SbRwhj0LhDDSRjJzo9oLeAc4JIIgrIEsggC54AijUebtiUb7pCQBZZIQKScGYLkCknDwd3a3UHr57JyS7Y5D7aNb+tEH4of3bKbnfPA9TecbX6PvM93ymGH/ctuq9ve5vjmsd5nW9fNG4o31zG8Hip8fneIyP/3z//8z//vdbdDURRFeXWoA+QthHJmBAD57W9/i4ODAwFA//u//8t/9Vd/5f/0pz/xarXii4sLds7RbDaji4sLLoqCnj17xsYYOjs7o/F4DGMMrVarLudj+CWPiIistWiaphdFAKCqqkvTmBlN01Auo4WiKNA0DYkIvPdUliXatu2HAFCWZX883bxunIhgrUXbtrT5hblbv5ueO2ZvFCq69YqiQBZ1bjrHNy6TYlfStrvxmxCRvhRWjLHPBemmN03T/S3dciIizjlZrVZwzknTNBBJZbCcc5K3IwAi5XJZIYTYtq0URRGXy2UsyzIaY6K1Nkwmk/iHP/xBxuNxfPr0adzd3e1FD/S/pd898QMAnZ6e0tHRES8WC/v11187Iiq996MY40REZt77uYjsNE0z995PQgiFpNJvivL6GXRq5XqEQIzp4T2kbYHVCvH8AnJ+DpyfQ7II0jlCOARESYHpUQRWAPIBJnhw28IEj+E76aVOxcH//R3Q65ul++mXl99of1ro7od+5zVeHa9K4PvuBJA3h1fZ5XqzANIteIeNvkIB5L7cRwC5/Xnd5na4Yr/bFrznc4q27Hv7lG3X9fqj6xwgNy+5ZvihfdPrhIYCCPCCAEJ0+bR0o4FzeStXIliHYG2qD8gMYQJMcn6ItYBNLg8qClBRAFUDFAXIOaAoIG0BLgpwFkIkJkFFRBCIknuEGYGTKB3QiR5pGLLgI11jhx3WKoQoN7DtM+4618W2aUPhY7hcN28zvH1zvzfN32zvdS6J22zjJq47zs22bC6/KcRstnc4/ypnxjZ3x6aotLlNvRlJURRFUa5HBZC3FFrnS3S3iRDSbyL64osvCAAODw/pt7/9LX344Yf46quvqK5rev78OQHARx99BAD405/+1AkDl741ee/7aZud+957dNtxzvXrzedzPHv2jJbLJRaLBZ49e9YLG845zGazfr1ueQCXpoUQaDqdAgBWq9UL3+Q6kSOEAACYTqc4Pz+/8RufMQbGGAJS6ayLi4sr15lMJgBw7TLj8bgf393dvXbZIXVdI4sVYGasVqtuunTzQwidW0TyvgQAOgFkuVxiNBrJ06dPcXZ2JgBQlmWs61q897K/vy/eewGAtm2FiOTZs2cyn89luVzKkydP5JNPPpHHjx/j5z//eS96AOvn1TsInZyc0Jdffmlms5kdj8duMpmUf/7zn0chhEmMcSYiM2PMjjFmpyzLubV2AqAEcL0FSFG+RwiDTsCu0yvGXAKrgaxWkOwAkfPz/LgAVqvkEgkhOdEklXKRGMEhZPFkCfIeJF3V+WvuOh8IIFeR3li23N39ssd9TbuG+x4O773fQTmh2+77una8dHtw+frfZd83LXfV/m4z7zbn5K7n4CbHw127eu57De67v6v2/aq6qG7frnUWz9Zj3zRk3Hr/t8kmSayPf1veyC2OgDbWGTg8blr7Vu8VGyLIcL2rnCZiLYJxiFWN4AoE55BT7oBcBmuYAULOIWYBhNsacA5UFkBRgKsK8B7wBaJrc6ksh+gDyBpEEURmkE3ltogIUSSV3soqdOcGiRh0hg7KY2nnqHJfrhMWriutdFPZpW1Oh+vW39z3bXjVNwpcJ1hct85N526bg2WbmHTVa1lf34qiKIpyMyqAvOUMOqy/i47re32bEhGcnp6+sO6nn34KAHj06BEBwN/+7d++sO7jx4/pb/7mb+60v88+++xW7fzkk0/w+eefEwDs7Fxd0WhTDLqKn/zkJwCAL774go6Pjy/N+93vfrd1Gx999JF88cUX/d8HBwf9+I9+9CP5zW9+0//dNE1/TY+Pj+Wzzz4DAPzP//wPAOAv/uIv5OnTpwIA//iP/yinp6cAgBxW/q4KGfeFAPBf//Vf8/n5efHHP/6xKsuyJqKZiMy99ztFUewWRbE7Go32dnd3d2az2awsy8rcVANNUb4nXrjzUKQPQEcIiE3O/zg/R+zFjySAyMVFEkBiTO6PEFLHWBSYEODbBqFZgdsWHCMol8K6bQfnNnItvRTie8Vd1rfZNnXHCkklv25Yt983KAUKb+ncvC3dvjnve1OIuYlOXY7E/flYz7tdq4YdsSy41bW5vO/t12Bz2av2u236Xa9H6pglhK3X4/ZXJ+0bYEhuw+3OQzr3qWTRXQ0j3fW/7f429y1Yvw7ipdewDP6/XVsutwswXduu2fdtrv9d2Dwnt7VIdsd/12uwfd/IQu3LCUrD96jr0ty2tdcbC28dQojwroE3yQFCnLI7wAzKmR5k7ToDpCwhTZOEkKpMTpC2TcOBCwRFAbIWxjkElxwkMRhEa2CMQSCGICJSEpUikigCQl8Si5A+N2I+T+oIUV6G6zrZb1vm6Tpe9XKvm7u4aG4zX0UORVEURXk5VABRruNe3zDzF7QX1r0pRFtE6Oc///md9rVNaNnGp59+2gsvN/Hw4cO7NIF+9KMfvTDx97///dZ9/f73v8cnn3zSn5vHjx/38370ox9JJ6p0PHr0CADwq1/9Cg8fPuxFDgD4l3/5F9l2rt+VsPJXycOHD2l3d9cYY5wxphSRMRFNAey0bbsrIgtjzGJnZ2f36Ohod29vb7FYLKaz2ayy1qoAorxREJDKXon0w+g90HpI0yYhpGkQVyvEZSp9JU0DNA0opAwQk8UTEoGPEU2MIEEvGBRC6Q7v+3Y05E5OD0LbdTx3dzXe5TiROjwNCVxcO1NuLNVDqbO9Ie473e+FCAwETiJc19F8l3OSO1dbIvh8HoC7dn0njAgsBO6214bSPfot0r5DviN8k7s6QGhwTm57PeTK63H355eR9Fy47fXoOrgbIoTBNbj9/iJsFDhEGMj9rj8YntP+By27vxtFBAZAgbgWQl/Yder43vYafBk68aO48/UH2o1rcFcxCsjXQ9Lr4M7XY6NNw9eHJ7r0hN/c6ubdRhGEIEDrfQpRCyG9voiyAEIA8zoA3djk6mjbJEaXJeJqCSpLyDINuxJZVBSXSmRx4RBzXkjMYkjI+SDRcBJAmBEAcL7uMYsdMQtGw1wUyOC5p52qiqIoiqIoynuACiDKG8M9XQvdOtf+gjs5OYF8N7cMbd3vb3/7263THz58eKkNv/zlL/vxXI5qc/n1ji7/SBUVOm4N/f3f/z0DMGdnZwUR1UQ0aZpmJ4Swa4zZI6K98Xi8t1gsFh9++OFid3d3PpvNxmVZWuecZoAobwSC1PkoSJ1cMhAxECOi94jtUABpEJsGaNvU6da2qVRWTJ2mMT+CAG13NzUxmASWCPwSb5np7vPU2dkywxPfWwBhibDZbWDkykI+l4gghE54YEak+72MSXIwfFzfbX8Xujvwfdf5n7Ol7lMSzEoSu4wIjHRbv54IIBCjYU53jL8CAYRFYEXA8VVcj7udh04MYwAm3PZ6UL4GjHZwDW6FSPqiTBEWdOfO9s790V1/T5w7nO8jgQ1fEwIbI4wQzBXFra57Db4MJAIrsb/+ckMpLOR2RKTz7/NzsWvjrfcLpOtBAGKE3QznuAfD14ffEIi2Odbk0ngSGkLwvbOiX59SDogw9yKIGIPYWrAr0nty04AKB16tIGUJWi5BzoGLMpXEcjkzpCxBZQlTFJDC5UcBk0WQEBhkOOWAECHKulRejALOpbGGWSciAma+XGJHhRBFURRFURTlHUYFEOVd4cZfwd+RdVhE5IUNbwodN7RFAHVufBeICD1+/Nj853/+pyWigohKAOOmaabMvLDW7o1Go33n3OHe3t7+/v7+7u7u7mw+n48mk0lJmdd9HIoypOsI5E5QyEHokkthifd9WSxp21RbPk+nGNbuEcG6A7H7+zuppqgoivKuIalcYBSAYy92CQhCuewdc8rpyA9Ym9x63oFaB25tEqmbBuQKsHOQImU5dS4QFCvQqAaKElymwPTYesBZiBnkjOTyW4G5L31FOZMktUsApt4ZIrJ2z3TiiL77K4qiKIqiKO8qKoAoykuieRtvJp348cUXX9jxeFycn5/XIjIWkan3fgHgYDQaPdjd3f1wf3//B4vF4nBnZ2dvOp1O6rouNPtDedMYFg3qit8NU6B4EKIZQwTFkKbFmASRmO7a5hBBuZwUS3dHP1BCUEqEk3Xexcu0lZDuFJcIWJKXK4GF7Dq45doMgUFEIYCJgNz3bTo7LqzEK7MWriPldghcFBAHxNjd+X+/0k82t+c2mPu2lQAAIABJREFUKQqEdB6sRCACgbbf5X2vEljyqq7HHc9DLv1k4+2vByE5Zly+ht01uPX+uut/D7dBf/0RQfl18CocIN01MIhXPheuew2+DJTfH2x+Ht76Ggyuf6S7H38n/Brc/3psbm/4+jBJNejnb9v6iyJBJ0Jfdoakcm+UHBrEaydICJDWg7wH2RbSGsC65AaxFmJdFj2K7AYpIEUBZEFEypwZUhYgZ2FywDpcDlrPbhPeEF6EGWIIkCzKYJ3LA6zLZVEWRtQRoiiKoiiKorxrqACiKMo7yenpKR0fH3OM0cUYS2ttFUIYtW07M8YsRGSvruvDxWLx4Ojo6IOdnZ398Xg8r6qqMMboe6PyRnI586DrfEz/cw7B5SgDR8cgUFOQQtAHHdhGBE4EpQgqERRZaDD36OzfhIG+o/Kq0jI3Hms3fk3Y81XrWhGQxPuLH/22bh/2va0dKacgwkaCIAK4X/d3F4J+l/PASB3/BoItZsUbW3FlEPorvR73OQ+3vx5dR3cRY86eiHfcn9z5vG/u2wlgEDauwf0zQIAcgn5Dm656Db4s3fW/7TVgAMjXPw6u/30yQF7memxrV/f6cLdozDbxY3N6JIIHgYmxEukdGKBcEssYIAbA++TgsC3gHcRYUBZD4FzKC8lCiKxWiM7lnBAHlCXgXApYdylgna0DrAFblwQPayAmuU7EpPD0VIqLEA364PdL5b26klhdeTEVQRRFURRFUZR3BO3kUxTlXYSOjo7Mcrl01trCe1/FGMciMp1MJnPn3G5RFId7e3sPdnd3D3d2dnan0+msrusRMxPRPQMDFOU7psv/oM6hQakzkogRITC5Ln1XA57zPdpdAC4JYAQ5RHgtfhSyDvo2uCFU6Zakzv/UUTms1X8fAWTb3zet290B/7I5AXfd97Z1N8Oa79Mi2hjedh0G8t3y2/d6HwHkPu14ndeD0TlB7r/v+z4HOhGEt5SYexkB5DZtuuo1+Cp4FdfgPgLIffd/1Ta718fdz872NYJQEqNZgJhdUtldIsK5ZGGABIZYixhNKl/IBtE0YGsRrYNYC3KuF0DgHFC4VBorB6KLTYHoVDiwdSDrkhvE2lQiy1qgyOHp0UKsQASIYhBMCk6PSM6PkM9BJAIjy4SdCDJ87qgooiiKoiiKoryFqACiKMq7Bj18+JA//vhjfv78ub24uKiaphl15a8mk8nObDbbn81mR4vF4sFisdgfj8fTqqpKa62+JypvDUSUckCIUkcnpXuiiVK5ldjVfieCEPfLGwAOhFIiSpF+aDvx41V0lA628V10XN52/6+9q+6KdrxJ5+BNasv7tu/vtE3XvAa/d17n6+AqNtr0ytqS6xMWkcEUU9kzQRZAYi+ERGL4GOCNRegyQthAjIWYVBILJrk7okvCBlkLuCR0UOGS0JFFD3LJLULZNYIildMiX0Cch5QFJEaIAEEEDIsggkAEcPociVnsiEjCkOTzlEpjpWOTTshTIURRFEVRFEV5i9DOPkVR3ilOTk7oZz/7Gf3Hf/yH3dvbK9q2rYhoRESTEMKsqqrd/f39ww8++ODD6XR6VNf1XlVVpZa9Ut4WaPORa7cDlOrMcxJCOIsfSQyhXgCxRCgB1ADqnPlhIbB4AzpKFUVR3mI6102BCCudcLCuNSVEkEjwxGgi5xB1TkIEMYTbVKqKGcKpbBV1WR/GgIxJ+SCuE0hSVkgnfHBVgooCXJagsgB8CZQlRCJEBBGUyiASoZUUnE5gBB6IQZSchL1vTASEdCzJeUiaE6IoiqIoiqK8VWiHn6Io7wIkIvjFL37BAMyvf/1rW9d1tVqtxgBmIYRF0zR7q9VqX0T2rbX74/F4N2d+jDmhv+SVt5ZLQkjv+sjxyPkGXwOsMz/QZX7glZa9UhRFeZ8ZitN9Ya2hq04IQkgB9mKSuJBF6v5922cxhBhkGEIG4DRO1gBswNaCjE1/GwdTFuDOCVI4cFkCVQUa1ZDRCNKMEKsWpmxhigLBuxSYbhhsDIwx8F0QOhMi8TojhDgJKPnzJeaSiiJaGktRFEVRFEV5O1ABRFGUtx06OTmh09NT/ru/+zuzWq1sCKEoy7JeLpdT7/1itVrtee/3QwgHTdPsxRjnzDyx1lbWWve6D0BRXoYXHCFY37k7zFy26DI/IsoYUXRB6HhFZa8URVHedwaltbZLAtLPkRggEBiJiBiK1tm9l6chO/lAlBwg2enH2RECNjDOpnk2lcqiogDqGjKZIM7mkNaD2gpoWlDhQFUJGANTOARjEIyFsQYehGg4l+VK5RMjxZQJAgzKY2UHSOcGUTFEURRFURRFeYNRAURRlHcBBmCNMXY8HjtjTLVcLier1WoeY9wLIRx47w+894fL5XJ/uVzOvPdFjNG87oYryn2gXKs9lZuX7P5AjjzPyyCLIDGCZS1+1DGgiBFWIsxgeUVRFOX7gbMgzTGJCkmspnW0Ol0e70WFLveJTZqUS2elaQzKwohYAxmNEaYzSOuBtgU1I1C5ApclYrMCO4fgHIxziM4hWAtjDIIxiNYicApzFzYIAGLeVYRAujJZMaZyi4Nj650hKoQoiqIoiqIobwgqgCiK8tZycnLCAPjbb7918/ncWWuL1WpVxRhHy+VyHkJYeO/3jDH74/H4gJkP5/P5bl3XU2YuiYhf9zEoyl3ohI/e4dHP2RZ4LOjydzk/bHZ9OESwih+KoiivBUJ6TyaJOWejk6zRly68vPRwGgHUAqCsMaznE3HaFBtI0wAhpFwo74GLixSOXlZAVSaHSFlAijIFqGf3CDsLsRac3SWBCUQMtgaRAM7OEOLsWskifCfaDHNCJH9mqRiiKIqiKIqivE5UAFEU5a3k5OSEv/zyS/OXf/mXtqqqwhhTnp+fj4wxo9VqNWvbdrdt230AB2VZHs5mswc7OzsPHjx4sLezszMry7JgZnWAKG83kkURDEquSAQkdkVW+uksAoMUeG5EtOyVoijK62BrmayN9+OXfXsmRgwBkOzIOL+AlAXIWkhdIdYjYDpBrGpIXUOy6CHW5XGHaAzEWoANYA3ImuQuMZyC2g0noYUIwkCMWQhhTvsdZFF1YeoqhCiKoiiKoiivAxVAFEV5GyEA/OGHHxprravrugwh1CGESdu2s+VyuQgh7GUBZM85t7e3t7f30Ucf7R8eHu5Mp9NxXdeFtVYdIMpbx3X9YsPyV939xCRJ/EjlsVT0UBRFefcRkG9B52ewwUOePwesBZgR6wo0mSGuVgiTCfxyieAcxNq+FJY3FpKniU1CCBUuOUWcBawFOQcxksQQ5CB3rN2JlAPTu7gQQRZjVARRFEVRFEVRvmdUAFEU5W2D/v3f/52//vprA6AAUC6Xy5H3fhJC2AGwALBnrd0viuKwKIqD/cTugwcPZvP5fDwajUpjjGFm/RWuvJ10JUcuTwSwTQRR0UNRFOW9QwTwHhIjIq9SKSwAoanR+ICVAE3TwtcVokuOj2gtonWI2QUiNosdRQEpHLgqQUUBLktQjIBzQIwQYxCZIWwgiBBmxJikEAEhxpiyqrDOCJHsYHzhM0oFEkVR3h5yHJ/g9PSUAODTTz9NlQzTe5l+CVcURXlDUAFEUZS3CXr48CF//vnn5sc//rG9uLgoLi4uahEZhxBm3vtFjPGAiA7KsjyYTCYP5vP54eHh4d7e3t7ObDabTCaTyjnnXveBKMq9EOnLp3T02bhpgfX04TIbfyuKoijvNiKCGDx8IAQQJLsw2hDRRGBJjLZt4ZdVCj7P4ekxuz/gHGBMFjwqUFkAdQ2qSrAPsF0pRVcgiKT1AUQyqfwWUXKBIK6zq0TW7kQiSJSUKQJcEj7UKaIoypuMiFAneBwfH9Pp6Sl9+eWXBACnp6dyfHwsJycnAoA+/fRTISIVQhRFUV4zKoAoivI2QABwcnJCR0dHvFgsTNu2hfe+ds6Nl8vlPMa4G0I4bNv2g6IoPqjr+sEHH3xw+PHHHx/u7u7OZrPZuK7r0hijZa9uiWhGxBtJF4SehJDuGqXxyyJI5whZ/1MZRFEU5f0gAGhASeggggchAAgCtG2L5tlz+FUDb21ybxiTylgZC+QyV+wKcFHA1DVsXQOjMXhcw4YkgHCIQBnBuXyWCJIYQoxAhAABd+HolESNKHmaJHdI72jsvnNsCiEb0xRFUV4jdHJyQo8ePaKf/exn9Mtf/pK//vprms1mfHR0RACwWCxkMpnE4+NjOTg4iI8ePZKTk5NOENEfV4qiKK8JFUAURXnT4YcPH9JPf/pTAsAAbNu25dOnT0chhGnbtrO2bRcxxj1jzEFZlg9Go9GD3d3dB/v7+3v7+/uLXPaqMMZYIlIB5A5QvoNTefPYfm1kY7ixDlQCURRFeV+IIMQsfrREaAH4KPCtz8MWgTvhI+d4sAFZC8plsFBW4LYFWg+0HhQ9SAQsgIkCCQFwDuwDorUgaxCYQcwgSkIMgFSCiwAmhkAgRCBK04SoFzku33yRP7FkUM5Rv5MoivL9QycnJ91vUT47O+Plcmk+/vhjZmbDzIaIDAB47+OTJ0/CYrEITdOEg4ODcHx8HP/93/89PHz4MKobRFEU5fWgAoiiKG8y9PDhQwJgAPB4PDaTyaRYLpe19366Wq3mIrJommbPGLNfFMXBeDw+nM/nD/b39w8Wi8XOfD6f5rJX5nUfzNsM5bs1lTeDS8LHNdel+4lFUPFDURTlfSMXpweIIAJEJEEihIgYIoQ8hHJ5LGYICMKcgs2NARcF0LRA8ECIKfcjuw0JAEIANSW4cJCiSCHp1gDGZMGDACYwJSEGzAAxwJTnCaQf574UVsyfXbLWP9Ie6bJA0o3pjRqKonwHUPd+84tf/IKPjo64KApzfn5ux+Oxubi4sDFGO51ObQjBLZdLBwDGmOCc8yLSNE3jmbmdz+c+hECPHj3yIqIiiKIoymtABRBFUd5U+Oc//zl/8MEHpixLu7u7a+bzuTs/P69jjBPv/SKEsB9C2Gua5qAoisO6rj/48MMPDx88eLC/kxiXZek07Fx55xHJd8gORA79aaUoivLewgAcIiAEA8AgOS4ISRxnAlgEDGTBQRAJkBgBpM8S9h5MDLNicHZ0AJLKV4UIWTWgqkwls4oS5CzIWrC1gGEQG4ihvrwWWZuEDjZJ9DCp9JYwA5zD0wEYSkNBcod0dWMkytAU0pfS2lY+S1EU5a50goeI9KWuPv/8c3r48CEj3ZBXlGXpQghFURRFWZZF0zQlgIqZy7yuX61WjbX2QkRWMcbleDxeFUWxAoBHjx55oH+LUxRFUb4nVABRFOVNg3LWhzk7O7NPnz51+/v7zjlXPH36tLLWjpummV1cXOyLyCGAg/F4fDAajQ739vYeHB4eHhwdHS1ms9m0qqrCOWdUAFHeWTbuhF3fT7YtDUR/aSmKorwvMNIPPQMBSwQhlZ7qarh0bpAIQUSaELNTowssZ0rpUSa7OEgEHCMQAsR7yHIJKRxQFOmRS2eRtSBjwDlYHcaArQGMBRkLMcllAmuSGJKXSSW4OAkh3ThR6ikctEto/RlHyB+FXbo6OsfL4BNPhRFFUW4BM3fvHfTDH/6wePLkCf/4xz+mJ0+e2KqqLIDKWls2TVMbY8oQQh1jrImo9t6P8mbaqqrOV6vVWVEUZwDOQggGAIwxAmCYCaIoiqJ8T6gAoijKmwKJCB49esRPnjzhxWJhARR1XZer1aqy1pbMPL64uJg2TbPjvd9n5sOiKA4nk8nBfD4/PDg4ONjb29vZ2dmZjMfj2lqrZa+U948+YpFemDwcKoqiKO8okoSO/ksQAYKIKCmDwyK5PiKloQCIEnJweRYcmAHvwciZUyKpBFaMgPcQ30JW2f3hsgjiXBJBrAFbC7EW0gkdNgWrk7G9UJLm5eWsSZ2PxiaxwxhEYyC8FkB6IYSSlCPIVpZc4ksgfcnOzdKdGqiuKMqQbaXzuveJnBlZVVVlqqpi55xr27YEUMUYaxEZN03TiR6jGONYRMYAYIxZNU1zxszfhhCctZZjjCCicH5+HgDE4+PjICKkpbAURVG+P1QAURTlTYBOTk7o8ePHPJlMzHw+t3/84x8La23tva+NMaOmacYxxmmMcd627cJ7v19V1YPRaHT4gx/84PDw8HB/b29vd7FYaNkr5T1Gkz4URVGUyxAAl9VxJwEBnZtiLYoHArwQGmJ4IYSYZ3i/zpESgZEI6gQQt+pFj/XQIjIDziEOXB5UuOQA6UWSJJTAuiSiWJfFkCSK9NsgSuPGIOTA9CSKJOEjxtQ4IUIciBydU2Qzv0xyJoqiKO8n24SPoXCaMVVVTWOMbrVauRhj2bZtJSIjAKPVajUhopH3fiwioxDCWERGRCTGmKVz7hkA5713lDfqnPNlWbY7Ozv+17/+NZ+enva3LCmKoijfPSqAKIryWhEROj09JQB8cXFhnj9/7gAUzFwx8zjGOHHOTUMI86IoFiGEhXNusVqtdquqOpzP5wcHBwcHh4eHu7u7u7OqqpxzzpImYr4URKShom8FV1yjbrJeQ0VRlPcezkNC7J0Tm71uQYAWBAtCEyM8CUQiIHltieAYgOBBrgVa27s6OidHJ2CIWT86sUP6oUvih3OAYbBzqURWUQCuAAoHcQ7iLKT1SQwxBmIjQi6L1ZXHipzLZKFzsaxFDyFcKYIAeR40QF1R3ieGzrDN3zob7wWGiOYASgCliNRFUYwATImo+2068t6PYoyjEMIohFABECI6F5G6bVtDRKZtW7HWhqZpVsaY5Z///Od2tVq1x8fHWb5VEURRFOX7QAUQRVFeCyJCAOj09JSPjo5otVrxV199VdR1XcYYq9VqNQ4hzEIIs7IsF+PxeHcymTxg5r0Y4+7FxcW8KIrFbDZb7O3tLRaLxXw6nY6YWbUP5R2Grhmny5P1ZaAoiqIAfTmsVBJre19bQPphSBLBURCYk0NEIiARiAzEkAQHn8pTxZzXISZleHSB5sKcylpxmp6EjgJkTQpJdw5iLNgYMBOMMTBlCVQ1pK5BZQkpkhiCokS0BjE7SyJ3pbEEngiRBZFTdgkxIYaQy2RlV0gcukIiiBmSytGknscc+j68YWB4hvQ7paK8uWwTN4H167ZzdQz/vuV2Xdu2+wAq7/3IWjspimJa1/VOVVUzIpp57+u2bWvvfRVjrLz3hfc+NE1ztlqtKu+9AcDOubharXxVVRd53mo6ndLnn39OG64TRVEU5TtEBRBFUb5v6OTkhB49ekRPnjzh3d1dBmDG47Gp67pcLpc1EY1DCNMY4473fnc0Gh3MZrMHR0dHH9d1fWCtXaxWq5qIxmVZjhaLxbiqKpfFD/0WqbxnUP+/PvkVRVGUF7hFpx8TwUBQIsJIEg4kZ2skAYQgMSASwTPDGwthghCnklRESfBgXgsjxAAzYBhiHdja9LdzIDYgIjgJsESwZQmZzhAnU2A0AqoKXFeQpgXKAtE7BGMRrUFgRjQGxlr4GBENIxIjRIBzZkhkymHp6W90uSBZ8OhKYTHQh6sTpbJa/WdpUoBecIrIcH6Hfv1UlO+dq3I8hsLCUPTYFEaG0zcygwrv/UEubzUpimJeVdXO4eHhwXw+3y3LchZCKLz3RQjBxRhd27ZmuVw2f/7zn5/94Q9/sOfn5+K9DyGEhpkvQggjESkAmKZp+Msvv+yqIKgDRFEU5XtABRBFUb4PCAA9fPiQfvrTn9Lx8TGfnZ3x06dPTVmW5uzszNZ1bUWk9t6PiWjqvZ9773ebptlj5gdVVX24s7Pzo/l8fpBLYVkicsxsy7J0RVEY1T5eju4OKWMMrLUwJgWSbv4oUN5k8h2tKoUoiqIod6BziRAEBl0nYp4hlHI2IsETgYgRg0fKCUYSDbpSVESpzBYzIgDigTvEmPS3ten7hghs26CAwFYlZLlCaFqg9UDTgr0HqhLiPaQoEJxDsAbGGHhjEEPoBZfIDBAhEMB5PFL6bsOUxRBOOSFEtO5xHN4dDkBi1zF6+XtP96kq/Wq0Fka6DtfhWvqdVFHuxVCc2Mzm2BQ3NtfZEDFemD78O2Yx9Ir1nIgcMvOEmWdlWS5Go9HefD5/sFgs9uu6ngGwIsLdo21bevbs2ZKI3J///Gc6Pz9vQgiN9/7CGPM8xliJiCMi473nTz75BF999dV3eSoVRVGUASqAKIryXUEAcHJyQsfHx/TkyRP+6quvzHg8Nl9//bXx3lsA9uLioogxFjHGAsAYwJiIZjHGnRjjbtu2e23bHoYQDq21h1VV7Y/H43lXQgsAqfPj1WGMQVmWGI/H8N6nTgbvEULofygobyKDp7/ku1dl4yUhg4eiKIqibNCJIDz8oJD8Xw5MZxBAETEm4SAAyXGRnRaCJDwIUhkqYtMLJMRJvGBjYQFYiXDtCjZG2IsCMQo4CmLbQsZjoG2ApgLKMueCOJBzEGaQtX15LWTHCRkGE/flsNgwKDtUJOeGJFMIp7ZROlJizh+ZlASVGNdOEMpGD1qHpw8dJRgui/Wncdx244h+VVWUSwzzODo2f9JdN284fShyXDXcJnZsrg8AIYRSRI7qup6Mx+P5bDbbXSwWu5PJ5HA0Gu2ORqMJcrySiBARwXsvAMy3334bjDErAKMYY52FjzKEUIiIRQpYp+l0SiqAKIqifH+oAKIoyiulCzU/Pj6mzz//nADw559/zgcHB/bw8NARkTs/Py+dc0XTNJWIVERUr1arWkQmMcapiExjjPMY4yLGuHN+fn6wXC73QggTALUxpnjdx/kuQkRwzmEymeDw8BBlWeLp06f49ttv0TQNmqZ53U1UXuCy8LEev2KoKIqiKNsYlom5YhHKZbKcCCBZ/MhOiCR+5E0BufwUgBBSx392jlB2lhoAFgLrWxgRUPAwxMnVsbyAvzhHXC0RqhpSFgjWIjqHmEPRo2F45vQ3p7JYyBkkyGIIjMnjaSh52Ikm6welZTqnCK2D1ZHzREApPH5YNgsECASE9bzu+HlwPjaFjxdctSqMKO8oN2V0dO7zzeWumnbTPjrXR/fopsVB6bttj+F2RAQhhIqZP66qarpYLOaHh4eLxWIxn0wms7Isx8xcbrn5LjKzZWYbY3QhBBdCcCLiYowuxmiJyBhjqCxLfdEriqJ8z6gAoijKK6ETPh49ekQ/+9nP6JtvvuEf/vCH3DQNr1Yra60tYoxljLEmotp7XxPRGMDIez+JMY5jjLMY45SZpwCmAGZ52o73fhZCKGOM5jUf6jsLM/cCSFEUKIoCzIymaRBCeN3NU65kmwiyRQxR+4eiKIrykjDSD0iGJNGj6zQcLJNMIxv9e50IElI5LUZ2nMQIggCtAOfPQW0DNA2kbdAGj7a6QCzKFHzuXApnzwJIF8Sehln8MGb9sCloHcYmx4i1IDdwjuTl1mJJyjHpxJvONXJJBKFURgucJI6UHxJzyLpsOWzq80aGOSMv5LLkrJEXUHFEeYvYzNu4royuiICZb8zr2LbtbdvqHjHGK4WNGGM/vxsH8MKwbduqLMsfWGvH0+l0vru7O9vZ2ZkURVEYY9x1ThQiYmY2zGyQymTZGKMREWZmatuWAODrr7/WF7eiKMr3iAogiqLcFRp8AaVHjx7Rw4cP8a//+q98fHxMZ2dnvFwuDTObi4sLY4wxZVm6pmkqIho1TTMmopH3fuy9n4YQJnk4LYpiNplMpnVdT40xEwCTEMJoNptNxuPx1DlXGGP4NR77O4+1FsyMoijgvcdyuYTNtbqVN4fhDzugS/7oZtLloeaBKIqiKK+IdZmsmyT1Fzv4e9tEHlA3HQAkILaCEAVeBB5AC6BtWsRiNRA6GGJSyavQBa53zg9jQcb24gdZC3auF0DIOVDhQDbNh80CSC6nJdktIoQc4p5KYnXCRz8dOWurK63VZYp0Akk/njJFpMsUyaWyokh2jwxCmYfneLPjd3N8mIGw0Sm8eU2GmSWK8rJsEyg2czqGy22Gjm8OY4xbRZLN/Qy3363TLbdN+Ohu3Opu7nLO9bmGnfAxFEO67XbbDCEUk8nkYHd3t57P59PRaDQZjUZlFjeufDExM5dlaefzeRlCqJbLZWGMscxsRIRDCPpCVBRFeU2oAKIoyk30WR4AcHx8TI8ePcLBwQF98803PJlM6NGjR/zhhx9SjNGcnZ0Za60NIbiqqiwAd3FxUcYYRyIyDiFMRWTivZ+EEKbe+2mMceq9n43H49lsNpsdHh5OR6PR2Fpbe+/Lsiyr2WxWjUajwhijDpDvkC4E3RgD51w/rkHobyZd6CqwKYJ0Q/2dpSiKorwiNspk3e8TRi4N0sZSOS0vQBsCvA9oVyu0zPCtX5e9IkpCCAHCWQzpSlsZzuKHhbABu+T4EOdAxoJcAS4cuCiyCJIFkOwMSULIuoTWWgCh9d9AygjpymTxQPzIOSJd+HsSR9YZI12KWve53YWoS5S0bH9WB53F/elZfwfrgtb74WZeAl4UQbaKJZuOExVIlA225XN0jo1u+lWh5MyX71cbiiWbw205HFdlenT76gSOTfFjKGwAQFVVqOsaOzs7qKqqb/9w+eHxDh7FZDJZTKfTcj6f11VVlcYYd935IiIqisLMZjP34MGDUV3Xo7Ozs3q5XBbee7NarQgAOefIGEMA8Ktf/UpfeIqiKN8TKoAoirKVHDKOLs8DAA4ODujXv/41ffzxxwyA6rrmtm0NAL64uDDL5dJWVWWXy2XBzIW1tlitViWAWkTGQ7Ejix+zEMI0hDCJMc6stfP5fD77+OOPZzs7O3Vd12UIwRhjrHPOTCYT65xTB4jyfnPFXXIiguGLg4aLa/UrRVEU5Q0lZYgQWmKsiNEA8N4jLldJAMkCRCRCoFSaKjIngYFoUMrKgowBWQcxJpW7sg5kHagokgOkTEPuRBDn0rrOAQMBBCY7PZiTMJJFj0gE0wkiWeRAHodZCycSCeDk/kilsbKQkrNEOkOMdFYQ0KXcEWyOD0ouPuRMAAAgAElEQVRpdZ3DPDh/a5FjLYKkfJINp01Xfms4xOCOexVC3jluyuG4avqmIDGcP3QiD0tdXbfutnZsK3+1rXzV5vTh352YEULohyEEGGPAzJjNZvjwww8xn89RFMULmSDbjkdEXFEUO845MxqNbFmWN/7+JCIURWHm83npnLPn5+fnz549G33zzTfFt99+a1erFTvn0LYtGWMwnU7p4cOHePTo0U2bVhRFUV4BKoAoigLkslanp6f0q1/9ih4+fIjHjx/Tr3/9azo+Pqavv/6aptMpPXnyhBeLBf/f//0fj8djFhEDwIQQrDHGElERQiiYuVytVjURVW3b1tbaUVEUs7qud4wxOwBmIYRJ0zQT7/2obdux9368t7c3OTg4mOzt7U3m83k5Go2ciFCHtZausx0r3w3q/HhzebHIFWUniL5MFEVRlLeUGIEQEGWVxA7KbgpO+RkRWRDoxAciIGeAsHV9WSvpHw7iHFAUQBZC2FkwE4gpCSFFASkKiE0uEnASVpLAwklKMAZM6+l95ggzxNA6hL2blh9gg8jrNqd1aV0mK7sxuvD4Tujoc0XyaUmOkXXeCJA7l6X7rtYJG2l5zmJL7/bI7hMRWZfR2hBV+mVVCHmruK5k1G2yNK5yYWw6Me6yzU33+GbZqm3jAHr3eVEUvYhx1fKbpa82BZDpdIq9vT3s7e31AshwX9sEnjzdWGsryjWvbvP7M7vouSxL55wzzrmSiIpnz56Z8/NzYmZoCSxFUZTXhwogivL+QsOyVqenp3R0dETHx8c0mUzom2++YQC0XC5pPB5z0zQ8mUz44uKC67rm58+f27ZtrbXWGmNs27ZlDjkvvfcjpHDzUQhhDGA6Go129vf39yaTya4xZhZjHHnvq7ZtqxBC2bZtNZ1O68ViUU+n02o8HruyLPU96g1BRZA3i6HEcfukDxVGFEVRlDcTAsAisMhlbAYiAIB11gYloT/lahAiAZSDy8kYCDcAW4jNIohJIgicQ7QWXJYpH8QwWAKcCMhaxLJEHI0gZZVKag1KYXWOEGQxo3N/pP11geumzxRJAglnR4mBmNDnlghLKqEVUymvLkekF3U6MYRyLgGQBA9g7SQZuDUkxnQ+0lnaqDC2/rs3iMSYRJxBia1L3/FyTkkvwihvNNuEj02XxG3K2G46PIbrDvdzlctj23auau+mgLEpRjjnUNc1ptMpyrKEtfbS/OF+NzM8hmHmzIzRaIS9vT1Mp1OMRiM4d20Vq0uHAuDWC3frMDOyWMIhBFMUBTvniJkp39R3x00qiqIorwrtXFSU9xARodPTUwLAR0dHBIB++MMf8ng8puVyyQCoaRouioKbpuEQAtd1zTFGk8te2RCCJSK3Wq0K55zz3lcAKgAjAOO2bacxxkkIYeqcm9d1vbdYLB4cHBzsV1U1Y+YihGBjjFZEjPfeFkVhy7K0o9HIadi5otwd/VmlKIqivG0QAIagkAiGgIRyLkhyf/TyPTMYqVxWPySCUM4DYANiBtjnclSmD0SX7AyJqwZkU4S7bRu4ZgW2BmE0RjudI9YjUFH02R+4JIZQzhghEOfwdOa0/b7kVirFJWadMRI7UcQYRE7lu8CMyAQRypkiKQelc4GACTGXuYqd8AFk90cX8bVRxqo7mQMXRy9kdMEhA5GFKe2DBtvut6O88dzGdTGcvm29zfyOq3I4bmKbM2RbhsdwOBQvhkKIMQaTyQSHh4eYTqeoqqoPLx/uY5jf0bEZqt6JKXVdQ2MkFUVR3m9UAFGU94STkxM+Pj6mg4MD+vzzz/kf/uEfzO9+9zsDwAAw4/HYnJ2dmaqq+Pnz5+bs7MyKCLdta0SEz87OTAjBiIjtHszsRKRg5kJEKiKqkfI+Jsw8dc5NR6PRdDqd7uzu7u7N5/OD6XS6W9f1xBhjRYRFhLohEbG1lowxt7IaK8p7Rx/sgRsNHaRyiKIoivKWwMgpGJKSK6IkAYSGwkDuuI/Z8RD7DvtUSgq58xPEIGawMSBisDUgbsDGwPgGhhk2Bth2Bbu6ABsLWjWQIAirBrEoIMYkwcNa0IbjgzpBxJicOZKyR2BtDle34DyU7A4RTiHrlEv6RELaHuVgaUpiTqR8/LQWKBiEmD/4kzbEySEDuiRqdK6OPmBdsBZOupJbyDoHMcDUC0vdcjGvH+nydwgVRd4cOtFiU6DYlpsBbBcKti0/FBm2bec6riuJNRxnZhRF0bs6Nl0rMUbMZjPMZjPs7OxgNpuhrusXhJqr2rbpVGFmGGPgnLvRnaIoiqK826gAoijvASLCjx8/5ouLCzOdTs2zZ8/s+fm5m81mxdnZWRFCcDFGx8zu4uLCnp+fuxCCa9vWxhhNjNF4722M0YQQLADrvXci4ojIEVGB5P6oANQARnVdT62109lsNjs4OJjv7+/vzmaznbquZ3VdV8yst+Eoyn3Z9htuQxDJP2chfS6IoiiKoryBdB2wAAylCG/JEd5GcnmovFiflYEcII71510nBoCyQyMQiBjkOXUYGwNeMYxhmBBg2wa2WSVxoG0hIQAXF0BZwuf8EBiLyJRFkCQUkLV9qHkngHS5I8jjYmzvPoHhfnpah5PoYdZ5IBFIwgphUOYL/ZC7yldZxODsBOmPl5JI0pe1ygKHIJcRY87DnJ3Sl/Ti3N4swjBfKruFPN67SpTXioiAeW2S7wSEoZui4yox46YSV8N1tgkZ25whV21ruA1mRlVVKMuyL2+1bZ3xeNyLH5PJBFVV3e0kvSU8ePBAnj9//rqboSiK8t6gAoiivOOcnJzw48ePGYCt69peXFw4731JRKX3fuScqwHU3vsSQNm2bSkipYgUItILIVkMsVkI6QQQA8DlZQsABYASSQgZT6fTyWw2mx8eHs4ODw8ndV3XRVE4LYD69rHtTjPlTYA2HnhBCFEURVGUt4VUDisV32fIWvzAZReCvPA/Ul2oziEpAX3xrPwdhk0WQgCQABw8OHiQEGh5AYoBWC0hrgTKCtG5VL6KuXdQoMsb4YGAkEWE3g3CnEUS7jNBkgvkcp6IdOPUlfIicM4E6QUeXueDpBNEvUBBgywPytsYLn8pJJ6SWAOThpLFGrJpXIyBuCTsBKRw+O68dvtTEeT1cl25quEywFr82BQxNte9zkGyLZ/jqmk3rR9jhHMOZVliMpngwYMHmE6nsNa+0JaiKFCWJUajUe8UeZvpnCidG6Vpmn7ew4cP9SWlKIryPfH2f6IoinIddHx8TIeHh+y9N0+fPnXe+7JpmlpERkQ06R4ARjHGmoiq7lEURVkURemcK4ioF0BCCCaEYEMIBoCNMdoYoxORTgxxk8mk3tnZGe3s7Ex3dnbG0+l05Jwz2fmh3bOK8pL0v1mvEDxEBLS120hRFEVR3lwIqT5rSuoYdNBesfzlJai3i1Cfk5Fnx7UfMokgAhIBosBIC44R4gOkCAghIGaRIGYHhSA7QXpHBfIwldyi3uFhQJzHicDGAEx9qatL7ouuNFVfqoqTjsOMSNSX3BJeOz6SWIJUxgrZOZLdHtK5YLr1s/MFnLJJyHV5JQ7kHOAsqCwgzvXiBwyBRNbrA2vxQ8PRXwubZa+2lb/qXCAhBBARrLUwxvQiw3Xbvimc/CpnyG3GgbUAMplM+vJWOzs7L5TC6o6xK1s1dLu8K3SOlt/85jc4PT19za1RFEV5f1ABRFHeYUQEp6en9NFHH5mzszO7t7dn//SnPxXMXBHRKIQwAzAXkTkRjYlojBRiXhPRyBhTjcfjejqdVs45hyR2mC4XJGeCdNkgJgeaWxExdV0Xi8Wi2t3dHU0mk7qqqkKdH4ryaklZp9vv7gPkmnmKoiiK8gYi8pJGRtk6eptVKATYGCExIEQPMS6FnudMDAFlF0dqofTltpKbg7LrgjhnkBClLHWiVKkKWJeiMpxLXtFaUKC1GCLMCIYRjAU5l8UIzhkgWZigQcks5j5AnUwSP5gYYINoOOeUWMC5lFFSlqDCg2IJAIiy3k40BqEbz9ekC6PXbxSvh+FPqE1RIMbYP7z3EBFYa2GtxWQyQVEUKIoCwNWlrja3dxd3x1Aw2XRzDOcVRYHZbIbFYoH5fI7pdIr081JRFEVRvntUAFGUd5yf/exnGI/HDMCcn587a23hva/ath0DmMUYFwAWMcYpgImITACMiGg8Ho9HBwcH4w8//HA8mUxKa60VEYoxcoyRRIQAcIxxGGbOMUa21pqqqsx8PndVVRnVPhTlu6PPRhcBqeFDURRFUe4FS4T1HiQCwx5NdnJ4YgTqhI91SSoiXgsHQA4X56RliMBKRCERtldZ1iHl3bArZzWcFo1BsA5tVaMtCohJpbVSI7lfLwkwqcRVJ8ZETu0Cp7JbZAzgbMolcQ5cFCDvgbYAxQhIhCFCZIJYA0jf2nX79IaKN4ZhDkgnVsQY0bYtYowIIcA5h9FohAcPHmA+n2M0Gl25rduMD/M/hvM3hY+hM2VTEDHGoKoqzGYzjEYjGKNxkIqiKMr3hwogivIOc3p6Sv/0T/9Ez5494xijISLrvXcA/n/2zqVHjuQ62+85EXmpW3dXcygNJQsjDATJ6Fl4IUA7Y7yYpbc9f8VL1vwM/wVya0CA8S2orWDBgAER9ix0wciakclh3+qWmRFxvkVmVmVlVfWFbLJv5yGzKysrMyLynnneOOckRJSiFDr6RLRDRDvMPLDWDqy1PWNMf2dnp7+/v9/b39/vDwaDJI5jAwAN8QMiQtXDLdUDABhjiJk5jmO21t4//2VFuQGoNS4i0JNLURRFUa4HEoFBAHkBQoCQRyBeeHug9rpAw2tj8bn05qjDeJngEYmHlYA6q0YtdAANEWSlEYTABs5GkDSDpGmZr6PyAAHVyc2xCHdVe6eUycwbyc2ZIXUy9irsVSgKkPdg7yASymIMgw0jOA+2DQ+Aqn1OpPQyaSTWVm6GZqeyWvzw3i8Eh1r82N3dxf7+Pvb399Hr9S4s9zyvkGbdF83XFkua1J4pF4Xlui88hHVUFEW5K6gAoij3mKdPn+Lly5fknKPxeMxRFBkAlogiAAkzd5xzPQB9Ihow804cx4MoigadTmewu7vbr/J39Pr9flwLIIqifHhWBA/thakoiqIo10+VF8QAAAUICIFMmXsDWM1/sXG88soAYCUgCgHWO1iEMt/IJQnGgGyE4BxQFGBrKtFjmSsEdY4TLkWPwAzHDF8lXhdmCBuINWXejziGxDHgHLgKmcQiZUgvy2VorDhePmOIlOG/UIbx2pR7Qnn/bEp+3vzNew/nHAAgiiJ0Oh3s7u5iOBwuwk1dRgBRrpd6PzUToCuKoig3hwoginLP+fOf/0xRFJG1lpiZjDGc57kFYJ1zMYAEQJ34vNPpdLq7u7u9/f39wWAw6A0GgzRNU2uM0S4sinLr0NNSURRFUd4HDJShqyTAAgjNhOpA6xZMS0GiwojAisAs/UUuDQUBO4eYMhjvIcZU4ajKP7IokKo8ILXwYUvPEWsR2CBUOT0QRRDnAFeAnKvEjwCBgJnAUQTYCJykgPfgIABXHS+IEETzit0UzeTnwDIEVv09hIA8z5GmKfr9Pj7++GPs7+/j8ePH6Pf7mmfjBmlHSFAURVFuDhVAFOUBYowR7z2MMXXs2NL73RjEcUz9fp93dnZMr9fjOI4RQvBFUUgIgY0xTBU3vR6K8rCh1qeiKIqiKNdFHcaKEGAF6zJGWwxpaQNUagjYEOTqEnULOARQkYOdq8JeteprNoUIhYngrQVFMcTGCMzwtQDiHMQZwEWlB4gEBAmlp4s1kPkcHEWQIgf5GCQBCAwyVEXaKj1gRETTjN0CajGqDn9VFAXSNEWSJHj06BF++MMfYm9vD3Ecq+fBLSGEQAConcReURRF+TCoAKIo95xPPvlEjDHh+++/D3meByLyjaEwxuTOuZyIMiLKjTF5Nb0gotx7L0VRsDHGxHFskySx1lqjAoii3CY2nY7UGhRFURRFuTQiCxGkmnDOvO+jbgF5gOEvnp0IYjw4RCABEKQMf0UEMQbBe4i3gA9ACAhAlficIZGFSRJQUUCcB4UyXBdDyvBXVXs0/8fNsSmvRi2C1AKIiCCKIvT7fQwGA/T7/ZtqrqIoiqLcOlQAUZT7jRwcHIT/+q//CkTkoijKi6KYM/M0hBADSEUkYmYmojyEUOR5np+cnOQhhCyKoo6IJCEE2+l0ksFg0Nnf3+90Oh1i7b6iKDdO/R4sUvdLJdU7FEVRFOUhUgkfCKEUOsps65CVfygfFYyB5DnYWvi8ABXV4B0QyjwoBJT5QKqcJiDSHGQ3RDvsVVv8cM6hKIpFMnQNVaYoiqIoq6gAoij3H3nz5o3vdDoujuPce28ATIuisCISV+KHEFEOIC+KYn52djafz+czEemGEFLnXLy7u9tzzhVpmgozhyqReh0+C83YpiJCVbxaKoun2t1XzbKKco3UwsdC/FAURVEU5YEipedICAAcJHDpASIMqUJeCaQUQKwBO4tQ5ECRg4syN4gJAeJLLxCIgAH42vsAUBHkBmmLGvX3OsG2tRbMvMgZotw89fuv9htUFEW5eVQAUZR7DBFhNBrJP//zP/s8z4ujoyPqdrs8n8/Ze09RFFGWZYGZHTPPRWTqnJt47ydnZ2fjEEI3z/OOcy4tiqJPRINut5uLSJplWQKARIRCCAyAQghc5xNhZjbGcKfTsXEcW/UYUZTrhCASsCJ66LuuoiiKojxcBCApPUAIAJMgEJXT6iTm5Q+QwkCMAUcR2DsE78DeleKHCEhQhryqDOrKzbPJq4OZ0el0YIzB3t4ednZ2EMcx9LXr5qnekQlY5P9QFEVRbhAVQBTlfiOj0QgHBwfhs88+83EcF0dHRyAiEpE6XmwAUACYM/NURKYhhAkzT0IIXWttGkLoFEXRnU6nvdevX/cnk0lqjElCCCaEYETEeO9N/d17b6Ioinq9XvTRRx91dnd3yVrL+gKlKNdBlWmVynBXdTiLxU/t04wAqYcP2UxFURRFUT4gZegqDqFMvk4AExBIyozsJIAniHOAK0DeAt4hOAd2pfghwZchtCoRZSX3RAigdjJ25YNARKXXLxFCvR9EkKbpYhgOh3j06BH6/T6iKLrpJistakFEREj3j6IoyodHBRBFuf/I4eFheP78OQDg7/7u72QymYCIgjEmiIgDkIcQ5gCmzDwlogkzj4mo65zrRFGUeu874/E49d53jDEJgNQ5F3nvIxGxzrkohGC999Z7H3U6nXRvby+NoigkSYIkSQBU72NVeKwKQPuuK8qVOfekWeQ+r80Uaq5QFEVRlPsMCUAQGBGYEGBIIERgksobpPLqCB5YiB3lIGEpftQSR50HhGrPA+3IdOM0c4AwM5IkwXA4xOPHjzEcDtHv99HtdmGtmnkURVEUpYneGRXlAUBEAiAcHh7iX/7lX+Qvf/kLkiQJcRyH+Xzu0zQtRCQLIcyJaCYiEwBdEUkBpACSEEI6m82S+XweV4nRk6IoYgBRCCH23seVGBI75+Jer9cF0Ds9PS06nU7BzF0RsSJijDEmjmMTRZE1xmh0LEW5BgTSEkVU/FAURVGUhwABYAgMBFYCIhAEXOZFBxaeIQgBIdS5QqqE6bJMes6oRBIJi3L1KeLmaYa/qr0/AMBai263i+FwiOFwuAiHpe9WtwcRoWauTEVRFOVmUAFEUR4O8vz58wAAX3zxhYvjWLIskyiKvPe+EJE8iqJZnueJMSYuiiI1xsQiEhtjYmaO8jyPnXORiMS16CEiiwFAUg2dEEIvy7Le6enpibV2MJlM+s65jogkaZqmOzs76d7eXoeZI6gHiKK8Pc2wV60zSaAyiKIoiqI8BBhAJKXkQaBKvOC1EJgElJE0q5BZFEKV96MSRqqy6uTnaHgdqBfIh6cZhqw5TkSLBOhxHCOOYw19dYthZoQQbroZiqIoDxYVQBTlYSHPnz8Pn332mQCQg4ODUBSFL4rCDYfD/OzszAKYViJHxMyWiCzKa0VkrbVxHNuiKCIAERHFIYSYiGIRSVB6inScc90oinpE1Ds9PR3M5/MBEQ2cc30A/cFgMCiKIqRpaqy1RERWw2EpyvXRFjtU/FAURVGU+w0BMJWoUflyIFT+oUFk8SwQGvNz9dTNVMWphZQpxmqhQwRUexNUidSVm6WZD0TzK95+aqFKURRFuVlUAFGUh4eMRiOgDIklw+FQvvjiC/+Xv/yF8zwvhsMhAzDGGNPpdPjs7MxEUWTyPLe9Xs8AML1ez4YQohBC5JyLjTERMydFUaQA0hBCB0APQG86nZ7OZrO+c26nKIodZt4pimKepmk+GAw8EfU6nU5irY2NMYb0Sf7WUu8afflVFEVRFEW5XZQCSCV9iCAgwFfGchEsPDmosQRJKX4s8n2gSh8m7bCaiqK8DXUIrBACWWvVC0RRFOWGUAFEUR4mgtIbhEajkRweHuL58+f005/+lF69esX9fp/G4zEDoCdPnvBsNuMQghERE0IwAAwR2el0Gg0GA+u9j6y1cRRFCRElWZZ1vPcTAJ08z7vOuV5RFGPn3BjAxBgzPT4+niVJknnvd3d2dgaDwWDAzAkRaReZW4jqUrcPWQtutS5MycapiqIoiqLcK5o5IgAYAiIAIqFKAkJVpjCBq2dCnTuEyoGwCJ1VeoFoxCtFeRea+T+IiLz32tdPURTlhlABRFEeNjIajTAajSAi8tVXXxGAcHBwQI8fP6avv/6ahsMhPX78mMfjMcdxTPP5nEMIxlprO52OYWbb7XYNM0fOuSiEEANI8zxPRSS11qbM3AkhjKthkmXZ+Pvvvx/neT6dz+cz772P4zi21kbqIqwoF7GM/9yWN6SSPERlD0VRFEV5sBAAKwIWD2YAQvAwCABCLX7U4a8WA1VhsJZCyGK+oM8VN41UIcjUgH43EBFiZmiIZ0VRlNuBCiCKogiw6OFfv92QiOA3v/kNDYdDevXqlX/8+PHCO2Rvb4//8pe/uH6/zyEEQ0QsIrbX65mTk5OImadJksR5nsfW2qQoijSO4zMROQshnIYQdiaTyWmWZRNmnsVx7LrdLrz3mbU2DSEYZuYoioy11hpjDKsyoigNloaIMmepAKA1dw/S7puKoiiK8uCohYwyE0jp9WGqIaB6XGgkPOfGMs3wV/oEcfM0Q9A2E6E3p6kocjsJIVDtBUJEFEURRIQmkwn97Gc/w3g81h2nKIrygVABRFGUTUhbEBmNRvT06dMAgH73u9/xZ5995n/729/yL37xCzo7O+Ner8dFUZgkSYy11sznc2uMiQBE3vu4KIpJHMeTLMsmIYSJc25aFMX87Ows7/V6Pk1TmU6nMyLqhhAia23S7XbTwWDQSZKEVABRlM0sX3ply3RFURRFUR4UjZweLI0B5QCUTw2LeQAgSMMDBHUwrEWR+lRxe6hFEFrkeFEPnbuA956YGXt7e/jb3/5GvV7vppukKIryYFABRFGUyyCj0UiePn1KAOSXv/xlAEC///3v6d///d/p888/x1//+tdF7pBOp0NZljGqzmbdbtd679MQQjeO40kIYSwiUyKaO+eyo6OjvCiKDMBpCKHvnOv0+/3+48ePd6y1bK01URTp9UpR1lg1R2wKfUWNQVEURVGUh8fC06MSQoDSg7ROek6yKoYQVoUQ0tCat5amh4hy+2BmMDPqXCCKoijKzaAGRUVRLg0RNZ+sBVWoLAD46quvwsHBAQHA7373O3ry5Al9++239Ktf/Ypev35trbUFM7ssywprbU5EhXOu8N7n4/E4z7JsHkI4894P8jzvD4fDnSiKsn6/H5g59953qnBbdXgsriJjqWeIolSsen3oi7CiKIqiKGV+sDoNOmOZM70pdDCw4jminSduJ+rhe7cIIVAIgWohBABNp1P66U9/ilevXt108xRFUR4MKoAoivIuSOMhfKu19dmzZ67f77s3b974brdbzGazQkQKZs5FZD6fz6fj8XjsnDsOIQxCCANjzF6n05kOBoO5c243SZK+cy5h5iSKorjf78fdbjeK41gFEOXBsy58SGNcURRFUZSHykLMECxEkMVv0vb2KIc6rJKGV7qdNJ/7muGwlNtJnQfEe0/GGOzu7uLVq1e6wxRFUT4gKoAoivLeOTw8DC9evPA//vGP8//93/9FFEUCwM9mM2eMyZh5Zq0dM/NJCGEgIgMAp/P5fPzq1auzN2/e7DHzbpZlO0mS9Hd2dnoi0o+iyMRxfNOrpyi3nOrF+IZboSiKoijKzUKCystDgIb4UbuEEKgcFfUCua00E5+r6HG7qYUPDVigKIpy86gAoijKe4eIZDQahSdPnvg4jvNerxdExCdJ4r33eRRFGYApEU2Lopgw89gYM82ybPb999/PiGgcQhgXRTHpdru7RVHspmnqO52ON8Z0TUkdDkvfBJQHhTSGiw5+PTkURVEU5WFRJkIXGAkwlUdHECBAVgSO5melk0CfHG4PzVwfzUFFkNtLI+yVoiiKcsOoAKIoygdhNBqF6lMODg5CFEV+Pp87ADkzZ2maTp1z806nMxORaVEUs/l8PnfOzbz3E+/9xDk3m81mc+993uv1XBzHPoQQut1ukiRJovlAlIfF+WGuaMu4oiiKoigPCBGwCGwIkOCBEOAqj48gUv5+w01UroZ6f9w96jwgiqIoys2gAoiiKB+SMBqN8OzZMzk6OpKf/OQnwXvvT05OnDHGxnHsvPc5gCyEkCVJkhHRjIgmxpgzAGMROZ1Op6fffffdaZ7nk/F4vP+DH/xguLe3x9baSF8GlIeF5vpQFEVRFGU7DMBKAHmBYYbxDnMJKFYSnpfPzwQARNpx4hbTfNchIs3RckdQ8UNRFOVmUQFEUZQPTfjyyy9pNBrJcDgMn376aXj9+nXY3d11aZr6oijcbDYr0jQtsiwriCi31s5FZEpEtXfI9Pj4eOa9d957l6YpxXHMxhi21lpjDBORhqZCAS4AACAASURBVMNSHiQaBktRFEVRlBoCYERAIkDwkBDAlddHaATBooYUImsiSB0YS7ktNBPUawew20dzn6j4oSiKcvOoAKIoyk0go9FIRIQAhF/+8pf+xYsXDCD84Ac/cG/evClOT0+LoiiKKIqyEMIMZY6QmXNumuf5dDweZ0VRBACh2+3aKIoMANPpdNIkSWJrLZG+DSgPjG1hrzSRqaIoiqI8UCpPD1ONBxEYEbjqZ8I5zwlSZxhrfio3SdPjQ0Nh3W50/yiKotweVABRFOXGICIBygf53/zmN+Hzzz93//M//xMAhCRJfJIkDkAeQshEZMbMUyKaisgcgBMRzOdzef36NXnv/Xw+948ePRoy88AYY/SBU7n3UHN0i1FCTwNFURRFUc5ltdsE1ZNIO1DcVvQ9R1EURVEujwogiqLcOJUQIiIiX331VTg4OPA//vGP3R/+8AfX7XZz7/1CAMmybB7HcTabzbxzTqpPP5vNiizLgjEmRFEEZkYURREzGwCs3iDKfWXVMCHL8fK0AomApQx3QSLbhRJFURRFUe4fVN75BYAHwRMhgLCeOqIRAqvxfTGqjw+3gk15PzQPiKIoiqKcjwogiqLcGmohpPoaDg8PwxdffOGGw6FLkiRPkiQLIThrrQOAyWRCzrkwHo/9bDbzANDv96nT6TAzS5qmvSRJEmaOoJ3XlPvKWuyKWvgov7IIbAiwwVciyA22VVEURVGUD8pC/CCCZ4YnRiAqu0w0n7xXoNVRjYB1o2wKe1X37VLxQ1EURVEuRgUQRVFuK/L8+XM5PDwMAPzOzo4AkOl0SgBQFAUzM6y1RRRFBREV8/ncv3nzxhNRPp/P58PhcJ+I9uM4NsYYzT73FuhL1e1mVdWT1m8CDgGxd4h8gagoENUiyIdspKIoiqIoN4YAcMzI2aAwBoVheCIILX8vh+Zf5bZTJ0FXJ3dFURRFuRgVQBRFuc3Iy5cvcXBw4L/++mv5yU9+Ir1eT05OTiSOY3jvxVrriqLwAFye5+Ho6MgXReGyLPPMjDiOk1r8YOY6FJa+KVyR+iVLuV3U+2S5b5r7SEAIMBIQhYAoeJgQNASWoiiKojwghMqwV0UtgrBBqMJgNeaCAAgi4Or74hdRQeS2oc/kiqIoinI1VABRFOU2I6PRSADQaDSS4XAYPv3003BychLiOPYi4rMsK9I09VmWuTzPfZ7nbjKZuBCCS5IEaZpGIhLSNO3FcZwaYywRmZteMUV5V1bCITSnN3pwlt/XB1UAFUVRFOVhIAACERwzCmY4ZgjV3SEE3HpmqD8FsgytKdWg3DgqfiiKoijK1VEBRFGUu4CMRiMAkGfPnuHTTz913377LZ2enmZERFEUMQCICBVFQQAwm81wdHRERES7u7vZ7u7uo52dnWGSJF1jjAogyh2mkfCDqGGQKJNi1iG6gwAOBGKGGINgLSLnEIUA1r6ciqIoivJgKH1CS9EjLKbVEkijgwQRpBEGS58WFEVRFEW5D6gAoijKXUEA4Msvvwyj0UgODg4ojuPMGCPOOYrjGM45Ymbx3ocsy8Lr16/DdDrFbDZzIoK4TAZiiYipAtoZXrlj1D3/iOqDtzyMy+lVQkyUBg4hgrCBNwZiLSACrodmzGjtTagoiqIo95JNnqArATMrbxARaUyXxYz6hKAoiqIoyl1HBRBFUe4aMhqN8OzZM5+mKebzOTqdDlX5QCTLsiAiPs9zP5/PZTabEREhTVPT6/ViZoaIBGttrOGwlDsL1aJH+bUdDkGqeQLKsBeBGMQMJoIhAgnBoIzzrQqgoiiKotxvatEjYFUAoZb4ISIgVTwURVEURblnqACiKMpdRL788svw7Nkz1CKI9z4kSeKJqIiiKBOR3Dnnvfcym83k+PhYjDGSZVmxs7OT9/v9vTiOu9ZaFUCUO0ctWiwMGiIgEVCoQmAJQJUoUnuCFCAQMcCMIIJYAAuBngCKoiiKcv9piyBA+TzBaHiBoAqNJcucYuoCoiiKoijKXUcFEEVR7ipSh8N68uSJxHHsZ7OZHwwGhTEmOz4+dt1uF957472no6MjTCYTmc1mUnmLxMYYy8x2GQ1LO8MrtxsClc4fdRgsYJn3o/YGCcuY3uWIwFfz5EQQYgiV0cBZ1AtEURRFUe4djTCXTeGjHupnBG783vYKaX5qqExFURRFUe4yfNMNUBRFeQdkNBqFb7/91vd6veKbb77JAMxms9mk2+2exXF8bK1945x7PR6P//b69etvj46Ovnvz5s3ro6Ojk9PT08lsNsuKonDee32zU+48zdBXbWOHJ4ID4AgomOBp1QiiKIqiKMr9QAB4AAUARwRHhECrzwUgrrxIGyIIUfW9CrPZ8AxRFEVRFEW5q6gHiKIod57RaBQA0Gg0kpcvX4ZPPvlEiGhGRBEzn3jvuSgKcs7h9PQ0YuZYRLpZlvHOzo7Z3d3tpGkaG2NUFFbuJG3DxEpvTqJFT1AhAoFgQAggVL4jH7StiqIoiqK8XwIAD0JBhJwYOREcCL7qJAGUnyRLL5Ayt1gZ+IqB8tmhTAwCAkH0eUFRFEVRlDuKGvsURbkvSCWEhDzP/fHxceG9nxVFcea9P2HmN0T0+uzs7NX//d///d8f/vCH//vTn/70/d/+9rfT6XSaOefCTa+AolyVttAhDe8PaXwvE6GXw3IeDXylKIqiKPcRAVAQYU6MGRvM2aAggq86P7TDYgGrnh5S/ZGGd4iiKIqiKMpdRT1AFEW5V4xGI3n27Fno9/vFN998k3W73YlzjoqiQAgB3vtkNpslALrOOWuMidI05RCCeO9DHMfWlKhArNxCtpggFj06q/wfRAhVL06pvT+qgQAYIhRUGkdIAEvLRKga51tRFEVR7hi0KmoUxCiIkXPp/VGHwqrDXwLlPZ+q5wcPACKL3GBAo5NF/fCgKIqiKIpyR1EBRFGU+4YcHh6GFy9e+OFwmEdRRG/evCFrLXnvKc/zTlEUnTzP+1EUJUmSJNZa65yTPM+xu7vb6fV6UAFkM6LG8Rtl4ekhy0AUVCc6pfJPO/9HvdxCAKligRcgZLU4IoCtfELUxqEoiqIod48y70cZ6iojRkZUiR9UeX9UzwbVzb4OdcVYPt+VzwpSPmdQXa4svEapegZRbgeLZ0BFURRFUc5FDXyKotw7iEh+85vfhE8//dRZa/M0TWdENAUwJqITZj5OkuR77/2ro6Oj13/+859f/fGPf3zzzTffnI7H46woCn/T63Db0ReuG2TRHbP6KlJ6e4ggQMqenCLLRKeV0aMeHMqkqHMizIgxo1II0YToiqIoinJ3CQAKlGGv5sTIiOFQdnpoPgcsE6Evnxvq8VoYAVWiCJXPfKVmos9+iqIoiqLcTVQAURTlXjIajeSXv/ylf/LkSeG9z0MIc+/91Fo7ttaeWGvfOOe+n06nr1+/fv3mzZs3x6enp+OiKPIQguYDUW4dtfeGLAwUDUMFc5nzo/YAaeT8qI0dngiBGYEZjsvQGBmVvUTzKklqnSBVGonTFUVRFEW5/Uh1Dy/v8aXXh1s8B5T5P+pwV20hxKP0DPF1+MyqzNDwDNFuErcH7YikKIqiKFdDBRBFUe4rQkTh3/7t33yapoW1NmPmmYiMrbXHURR9b4x5nef56/F4/Ho6nR7neX4WQlABRLm11CGwQtNAwVRNL0UQMJfiB7BIeO5rMYTK0Bi+CodRECMnRk4GGRlkVcxwDzVzKIqiKMpdYZH/ow5zSQxHXOX9oMVzgUfZyUGa06vvAYAwl5+NUJtAGR5Tk6EriqIoinJXUQFEUZR7zWg0Ci9fvgwnJycuSZJ8b29vure3d9bv94/iOH4TRdGbKIqOoyg6s9bOjDEFEakAotxOqlBXi2SnIhBZzflRh72qjRiL8aZXSC2GEKFgQsaMGTPmbJATlwaSm1xPRVEURVGuhKD2BG3c61GLH0vhox7Q6CyxGIDyGaORVL3OC6JeB4qiKIqi3FU0CbqiKA+BcHp66j/66CNnrc1EZMrM1nsfF0XRdc71jDE7AE6zLBtnWdaNoii21hpmNsz8YMViIlq88Nafmvzy5liEwZLSEFEbMKjy/IAxgLUgayHGgKpx+ADxvhJLaOEpUk4QhBAQgiCIX0m0riiKoijKHYFQ3r+NgTADVD2+chXWsn5OMLb6LJ8TwFzOw7zoYEGEMgk6AVXQzfL5QJ8NFEVRFEW5gzxYo55yLdA1DYryXhmNRnJwcOCPj49dCCEnovnOzs44iqIzY8xpFEUnIYSTPM9PJpPJ8enp6enZ2dk4z/MshKAJ0aGxhm8DpSBR7Qeq0pESN4waDI6ilYHqwVqwjcBxXBo76sGUA7Mpi6lrENGLs6IoiqLcJYhKIcMYsC3v/xxXzwRxXD0bxIvOEWQtyBiwtSBjQcyLnGJgrvKOlZ6lAFT8UBRFURTlzqIeIA+T67BrqW3sw6NvHW+PvHz5Uj7//HM/Ho+dcy4TEXjvY2PMiYh08zzvHh8fp3/84x+7w+EQw+EwfPzxx8O9vT1jrY1uegUUhYiWV4FKCxEAXPXo5CgG4hiUJCDnQIUDB0GovD5ABPa+NHh4DxYBB4H1HjEEHS9IJCCSAAMVQBRFURTlLkFEIGMXQoepHZgrYYSYEayFRBEoTcohScFJApPEMPFSHJG2lymgAoiivAUiQiEEfaxWFEW5YVQAuV8sbqzN0CVfffUV/f73vycA+Oyzz+jzzz/H119//VY34eFw+N5u3p9++umVn6p/97vfvY+m3Dp+/vOfL7bNq1evVrbT8+fPAQCfffaZAMDTp0+rCDbLw+GDNPKW8/TpU3n+/Ll89913/he/+EXx+vVrcs7NvPeTOI5PQwjd6XTamc/nvaIoIhGJ9/b2Uu9996bbrigAFiEpAJTiRwCIGcIMNqb09EgSoChKgcM7iAhClTMEzKAQQM6BQ4AJAisBtnCwhhERYI2BCWGZAeSKV/x3udg8hDfD9xVWjDaMAe39cfW6L7dPHsKeuy6ua/9fxza/qC23db/KhrF16BLzKMpdpXl2LvtFEGAjUJzAJCmMjcpQmACYCUyEYAykEkAQx6A0BXVSUJLCJAlMHFfeIAaocofVn3X+MRVBFEVRFEW5i6gAcj8gABiNRguh4/nz53j8+DF9/fXXdHBwQPv7+zQYDAgAXr16RcPhEADQ6XRW3nCPjo4IAM7OztbefB8/foxtv70rg8FA/vCHP1x5ueFwiFevXl13czAYDFae7ofD4ZWe9v/6179eeZnzePXqFR4/fixAuR9ms9mi7H/8x3/Exx9/LABwdHQkL168EAB49uyZvHz5UgDQ06dP5aELIkQkAMJoNPLee3jvEUKYM/PEGHM2m806IYQkz/OOMSbpdDrdoij2RERDYCm3h0VuDlrmAmEu837EEbiIgTQBeQ+EUNop6njg1pbih/cwIuAQYEVgiwK2iGCsgak8Q2rknQSQ22JAfddL3sXr0Z5jc42yFEDOKXL9p/PrXzGENcOkrbXjatuBLr3EbdnPd4HGFr3qZlvbGbSxmMvts8seC7dx324/qhf5qprT1pbYWMwN0GrApTb1Ne2PD7H7b3r7bmq7nPv13Yr/gKcKyaqY3nQMhS09P2yaIlQhrZgIgUpv0cAMRNFCAEESgzodULdTiiFxDI5joMohQlU4rEVusBBufNcqyl1FREi9QRRFUW4OFUDuNgvh4+DggF6+fElffPEFDYdD6vf7lCQJ/+hHP6LZbMaffPIJZVnGk8mEiqKgKIoIAIqioJ2dHcxmMwKANE2p3++j3++v3Jjn8zklSQIAqD8BIMuyK93AkyTZ+tycpumVn6knkwmePHly1cUupG7LeDyuJ620rdPpyOnp6dblP/nkk3N/vyzdblcA4OTkBMfHxwIA/X5foihCURRS1/X69WvM53MZDAby6tWr8PjxY/nuu+/k4OBAjo6O5Pnz52E0GgkAjEajtfV5QAiA8Nvf/hYHBwcym82yEMIsjuNxCCHN8zwhop61th9F0Z61NmNmFUCUW0HT4EGE0qBRhagQZlAcA86BpYzWzVUccLEREEdAloODB/sADmHFC4SdB7xD8AFlP1IqbzB0jl1nQ16YdxVA3l/i9bcvlzatx7ZVky21LaKHhAvFj23bsD3W/N5w/9zSONnQrov31mLauTmAWl4nH6B38Ifwf7j+ujcZvLe3YtMvtJi4TKF2mfaslyVbKrhwwpW5tvxRsjaC9tHerIu2zFNOWz1R35/n2rqRuu2jJRcXcs6eppX1vHh/tdd785rT2siG386duvn4ak+6vivFeQ1t+UqsVLptC7xLfdfP2tYVaVwLltd2QhniyhiLyBqADQwRPIBAhMBLDxBEESQuw2YiTUDdDiTtAGkKiiLA2nIZokX+j1oEIXyY67yiKIqiKMp1ogLI3WPF2+Ozzz6jJ0+e0Hfffcc7OzsLwQMA/+1vf+OiKBiAmUwm7L1nZuY0TckYQ3mek4jQ2dkZGWMIAIwxlGUZOecWz9tFUVCSJCiKAs45iuN40RhrLZrzNmkKJTXe+41PzCEEKYpi60pHUbRxuTRNJcuyrcu9LSEEAQBjDABAGk/6URTJ2dkZiAhxHAsAzOfzleUnkwnSNJX29KsQx7GcnZ0t6q8Fj+l0KkmSyGw2g/denHMSRZF0Op1QFIUURRFevXoVer1emM/nAYBMJpNwcHAQjo6O5NmzZ+Hly5fyUL1CRqNREBH56quvws7OTt7r9WbGmCiKoth7H1lrU2buMfOu9/4sy7K5tTY3xnDF0vKkKDcBEUIIlfgByMIDJC7zehCVIbGMAdkIFMegLAXlOciXHiAcBCwCEwQGgAkCCmGtnrYBnIgWVvo6OeoFjb3E+lSf7y3x+iZj3Eq/8Y3tWV72N5gfNwlDAkBko8F1uYxc0ti5/q00Oq22SBbbbP1vc6w2kbWNryvfNmx/Wv2ztcXtbbNiHLuKof2SB8CVjpMNhvMrsa2tLWeOTRLTloY0yjz/eGjZapf7VzYJc9ScdWs55b65ggvAeRv7YoemFVHinR80pFlp2/jfqLM13pYhFtMWRV18RJXzrK/BxUuuHhlvI4BsFjabRwBt93TZWt52tgoglzR6r+SrekfeWkDbdN3aKBq8Pe3r3lWXPk9EaF+P18YbB3C97wWAAVDn7GAQPJUJzAMRPHPlDboMg0VpglCJIKHbATod+KgMnSV16Ku6/Lq9Kn4oiqIoinIHUQHkblA+64rgq6++IgD85MmT2gjLANgYw/v7+3x6emo6nQ6/fv3apGnKAExRFNZ7z0RkkiThLMs4hMDWWs7znJiZ0jQlAGBm8t5TCIEqQy/qz7otGx7YVx77o6jMF10UBRljVma21m4TOs59mq4FiTbOOQlto90lsNaulddqlwClu7iIiHMOAGCMkTzP4b1frEsIQTa9oOV5LlwnH7wC9brmeV6HbQIzCwCp6pQsy6SeV0TEGOOLohBjTAgheOdc6HQ63lobvPchhODn83mI49gDoCdPnsiLFy/koYbJqrar/Ou//qv7+OOPsyzLpkdHR7G1NnLOdQAMnHPHk8nkNI7jsYj00zSN4ziOmNncdPuVh0kd8qoeBwAhAQwDYkpjBkqvEGMt2BhwHIOyBJTnMEWxyP9BIZRhsARgAQyoHK/KLstpmNgIICqvZ8Tb7R+lIeZqlqDm5ZM2mHxErn6NX2W91++GVmwcbQoOq8auDaJIXazIar/ipqBSW64usPdTbbxbaSotev2W7Wk2dL3NTTv9ZhP0Bb2/m+Ote1xbYlkTT7ZZpts1tLf1exVA3oFNFa4JIJcUP1ZEj6sKIPVOpbV90BxfPWwae39xcDRbu+042Lyfti12CZ2kas5lJYPtE9utp3a5svnY3bSPrmLLvbotflvhG6Y3jonNhvH2Pt8ugF3YqksLGecWsmH+LdckbB5/V7YdSyui0sY4jucI1Vepf+uXy5V94W4gAI3XH2p9SuP9pxYopCqYUd7PPUoBRLj0FPXMCwEkRBaIY0gUIaRJOSSlIBKMgRADlZdpkOXZc69fEBRFURRFubeoAHK7IWDp7fHVV1/RkydP6lBW/PjxY+O9Z++9sdaa2WxmmNkws0nT1AIwzjnrvbdEZKrvxhjDImJCCEylRYuyLKNa/BARBoA6PiUzU5ZlZK0FES3CXllr0Y5hSUSU5/niu/dl9KDKgA8RkXpa/b0ed86hLZg0f6vLaFIUBYwxC4HismwSVJr116JK3T5mXhFBACDLMmmu13nlvU3b6jJr7xjnnBhjasFDQgjinAvMHJxzIYoiXxRFAOCLovAhBC8iPoRQj7udnR1/dnYWTk9Pw3/+538Ga204ODiQ//f//t8iTFYVIgt4AO84w+EwZFnmiqLIAEy991ZEOvP5/Pjo6Oj7EMKrs7Oznd3d3eijjz7a2dvb61lrzbWF9FCUK7LI+1EZJBiV4GBMOcaV90dkYaIIpijASQ5TOFBRVN4fofQUCQFGqDSUVOIHL8SPhoG/1ZO29PyQhQfI6tVvgwF203o0RtYMuRst4e96OTp/+ba3x3J0kySzXKbdyXi9w/QGIaQpEW24lKyUuRA8KvFrYdhtbrWmgbsxZeNl6nxT5EqYtWrYtDs2yD/nrtOy7HMMlvXiW6+vy97OV+L8PhsXs1Hl2lTuRRVvE0GadW2RJRoWXZLm1m8a91cLXOnsvlUEuL7b/IoI0Sr2qrUszkZqH9v19AuO5JV5m55qGyQQubiNy3ZcZU2uIH4AFwog64JX+7M9fl7TLg79tP0aUl8XLi+AtCdd11F33rOYtHbZpnnfpR1rpS3qu3ypsuUyUJfX3M6Lvb1yS5FFdbXwIagED5GF+FF6gJReILUHSFiIIBF8JYb4JC7DYlkLMVyGzKrKvvcvBIqiKIqi3HtUALmdEAA6PDyk4XDIBwcH9Mknn3Ce52ytNdPp1MRxbJjZhBBsnudWRGyn0zF5ntsQQhRCsMYYG0Kw9TgAIyKWmTmEYJiZRYSNMUxEFEIgKt8QuPJ8oOb0WrioRY/KQ2Hx7F5Pr8NGtSmrW74ZNMfbQsmmZZvzXfa3lY1KtFJ2u65NbWgKIM3f29ObAkm73E3iyHnU5TUFkHrcWhvqMkMIEsofvTHG53nuRWQxMLPLsswzs2NmVxSFOzk5cSEE3+/3vffe93o9n+d5+Id/+IcAwP/qV7+qc4WEp0+fBgC1V8i9fPd5+fKlHBwceO99HkXRbDqdWiI6m0wmJ0VR9M/Ozl6fnp7uPnr0KLXWchRF1lprK6GRKg8fVUOUD0pt0CMAQgQYggQBcQQYg8AOxlpQ5EuPjzguk5sXDlQlQKfgwQGlEAKAUYbLIJT5P8r/tDQaUduAJADRijGmaTrfYopdXY/lCq0ac29AANnWm74pVrQv5Svmxy3GrxVDYTVPfdVoGxhXDF0NQ3LT8FVvqaaYsPq32ebNPZ/Pm0aNdSj3f0u4WP3YMrZib99gKN0Q+qW5Magh+JzXzquwQaS7NNcigGwYX2vGcmevnQGLxetzbnmO1Z5ZTTPpSm0r6tK29l0fK4Jc9Wf9bN5Q9wYhUWR53Vk9ple3J6HWeTYLMOe2t1JTLpBI378Isrj8bfGhW9uR7bnOO65bbT/P8H5OkVeSWs7ZTJepe+HleEHhW71ALrG7rvXh7ZxrY3u2FcG9nLBxxvb2XhXBy89lf67lQcyQRQeJ+khhLvN5CBuILT1BgrWANYCxZc6P2IJsBFhTCiBECCB4kYV3SS20vIU7lKIoiqIoyo2iAsjtggDQP/3TP/HPf/5z+tGPfmQeP35sj46OTFEUNkkSe3x8HMdxbAFE3vvIOReJSOyci5xzEQA7m80iIooqscMCsMxsRcQSkQkhGBFZCCAAmLYgIsTMqIUQABBZ+pPXvzdp/r6yckRSixAhhLYgsfUVpS1cNENeNX87LxRWs95t5W6al4ikKX4ApcBBRBJCWIgV9ee2Mra1a1ub620VQoCUSpSEEGCMCUQk3nsQUSiLKEUQEfFEVH+60tnGO2YujDGFMabw3jtjTBFFUeGccyJSeO9dmqYOQHF0dOR+9rOf+d3dXffrX//af/PNN6GVM+ReCSGj0UiePXvmDw4O5L//+79NHMdmNpulRVGczmaznnPu+8lksptlWdrpdKwpXXBMt9uNkiSxRKTeIMrNUBlM6t6ebBi+MkpYZoQg5fXHWlAUwTsHpAL2HiEISAIQaqMGAVWi0/oq1jQ6LsZ5aZBqaxQLc85lwttsFBJKM822nsWrtVw/G41WG0MHNY2z0p6tIR6s0g6J1RY/mstuCjdFQovewqWBdIPxc2FIo4ao1Cz+cv2vl3W09ufK6Pq2aQo3q5tkXQBpf5XWuq8dRS1B5d2uuu+y9HUIIHUzthlxt/TObwhgK+NlCSvn4MaaV4z870n8aB0jzbqbSHvill2yPCxoIaY0l2+KEkuT8vbcRGtHItGFHfaX2/MSj6yy9ctqmc3fzxULV6evnh1vI4Cc366LuKYz54qVbqt1uwiy7fy5djY0rXkdBDbf71bvn5s99toehovrckvdXDsvFkLF0htk4cXBhEAMqcNgVTlBvGF4U3qF+CpM1or4gVJmFAkqfiiKoiiKcmdRAeT2QIeHhzwcDrkWPrrdrnXOJQAiIkqzLEviOO5471MRSQEk3vukKIpERGLvfVwJH4uBiEwtfIiIERGDsgOqQenpQdUnqpBYzV7ti7es2iOk/qwb3RY72r8vVq4ynLe9IbZ5R2wytG8SC0qN5lJvNWszbaqjKqvdxrV5G94ZdRtWfm/Of9l12VR+LXzUdTSFEWDl3cYTUagFEGZ2IuIBOCIqjDF5JYTk3vuciHJrbZbneWaMya218/l8njnnsn6/n81msxxA3ul03GQy8U+ePPGNEFmLTmD3AHn58qUcHh6Gb7/91k0mExfHcea9n4UQJsaYU+/90WQy6X733XdRHtePSgAAIABJREFUnuc8nU7p0aNH/f39/Q4zszFG3wSVD0/ZNR+oQmL5EFCL0VQl6w3AIg64YYYJAWQMWAS0GJYXe5Iy70dbDqAqoSpo2aNb0DKCvKVBZNWY3Y5xf3GYlvUCt365/HIXrMqqF8Z6Aat9s2tTZ8sItsGGSa0ZFkZPWRU96r/LLdQ2ttG5u2OzMLLsbrxiVl/0qJd2A5fT1yrYHjZspb4NMyx6fW/wEGkLT9vKv5gPIYCc9+Oq4X8pXFy+6nK8cZQRbzfPrxzbtGmOd2ZFIFhZvdXwU5uadW4Yo5XFluF+6mtcu1RpqDwr4bMa86wJGpfQMta8385t8GVoHQMbBNZNtK7Ml63sysgWI/fb1tgUp1anXH7Zt6mvybok/A60xQps2n+06eK3aItU11TaMC8tZ22JioAEacyz4exq5eqoXxSEyk9wJYAwITAvBm8YjgmeCQUBDoCX0pMkAFUOkLe4JyuKoiiKotwSVAC5eWg0GhEqO9XBwYHJ8zyaTCYxMydRFKXOuQ4zd51zXe99H0BPRLoi0jXGdIwxnRBCIiKxiEQhhBjAIvxVLX4A4BBCbQ+rvT/qsFd1snOqQl+tiBn1ZzPnR1PoqF8OK8P82luGbLMUbWajqEGbe1RtTEC+YdkL6zynMWu/l70GRapttDV017a6z2tzQ+CoPVAAQGrPk3p6Q3gJzBzqTyLyTSGEiApmzq21mYjkADIAM+/9nIhmAGZENPXeT4loOp1OZ1EUzUIIMxHJoygq8jx3/X7fP3nyZOERcl+EkKdPnwoAvH79OkynUxfHcc7M8yRJJnmen4nI8Xw+73z33XfReDw28/ncRlFker1eVOXaUZQbQQBQ3TuTCE4EppoeiOCZQSjzedQ5P6gKiwEJK+IHqrLaRqKF98ciHMnSlLVsxzYT58W0hQJqTX0rc8uKjfr85Zv1yZqR/+JlVmZvLH/RerR7/G4TP5q/yWJ/LUvfvHa0xfa2NJy1m72xLdSoq2WkbZfSeBhYqW/T5myH1GrWt1LuStKHi9fj8lyTALLh67aaNpr+W8LPujn/guqbm2clDNaGOqUtCLyfW3dTX2noFisNadd8WQGkFjea4sdGb5cNz4/NcqjKYXSpui859aqzLGbcUP2K1NI657acddfOtlW4PgHkvFou15Yml/IAuXyVl6hwdXz9Wkcbp2+6dlOjjLW7C60KHa1qz/UYEloKIM0BVVJzoVoEKccDEzwRPErxIwDwaHqTVOMi5543iqIoiqIotxU13t0gIkLPnz/nly9fmp2dHbO7u2tPT08j730SQkjyPO9473shhJ5zrh9C6DvnBiLSJ6K+tbbf7XZ7vV6vx8ypiMR1/g8RsSEEC4C99wYNwUNEuBIvuDLkL0SPCqp7/NYiR92z+Dzvj8uGPrlMGKWL5rnIg+KybPDsuHCZtiDS9kLZInisTLts+9ueJE3PkEa9UoXDEiIKzOybQggROWttISKZ934+mUxms9lsmuf5NIQwjaJoEkIYM/MkhDCJomhcFMU0TdPIWjsPIeSDwaAYj8dF7RECIDx79swfHh6Gux4Wq96Of/7zn0On0/FxHBdRFGVFUcziOD7z3p9kWdaZTqdxnudRkiSd2WzWCSF0cQ8EIOUOUydEx9K44VH12qzyczAzKAQwl9f0StFGmfGjYWgRKadQu4p26BlZFUNkdd7Lcv61dt1IduUTrWF9vdiYR+0J57IibrSFClqfczF66dBeG8QBVMazZuz4cwWb7YnQVw1n68pHs6nU3DStAldFms0NWdS1qnKsztMod034Wd/M7ebeas4VQJrzbRFAmvuJNqoLi1+3ix+tiauiwfu6hbW9NRrTN8y99DRql7IcWd8+srouG+fB2ua6jNjUFlYuzZUWWhfC6q9bxcbLeTy/A+dfC99VAFnfPpd45j7nt233nPb+vmRVl6aZG6p9jVq/BTTy9aDp+dHa1g0BpCx/7Q61RRDZvA1CyzukFj+wEEYIgVAKIQQIl+JHHfoqyDKZ+oqHi4ofiqIoiqLcUVQAuSFEhF68eGEmk4n9yU9+EolIxMzxfD5PmTn13ne99/0QwkBEBkVR9IuiGIQQdkSkz8yDNE0Hw+Fw54c//OFOt9tNjTFRCMFUA1deH1SN1yIH1eNAbQtb9+RAJYK0f9+2LhuW3zr7lTfWe+Sqxvum58mGaddSxznLSXt6WxCpPEYCgPozEFEwxrg8z/PpdDr77rvvxnmen02n02kIYeK9nzLzGTOPmXkcQhjHcXw2n8+7URRNrbUzZs4AzAEUcRwXBwcHxWQycS9evHCj0SiMRqPrUaRuCCKS0WgUoihyIlKISMbMU2vt6Xw+7xpj4qIoYudcKiI7zJwRkcctO56VB0jDW8CjvKjXxjtiKj0+jCnNo7Q0r5Q3gEo6qcKdbLx6N4yHdc9pqpIGr814vSv2dr3UpTl68fIrBqQr2XVWjVNbQ9hcwiNic/VL9aNt7Fray6rpLY+Rc5p6rsGs2St5MVfTgn/O9jmv3HXL4NqaViOb12ODffBWc1ET18OhLQ20mzyFFmHNuM5X0Z6nPqvPrbSubMPE66aSF9oizUV26M3KSEN83TyTrM5QLUZbp5/bhnfhbcQP4MIDZlO+nQ9CHWbxWoq64Br1DuXWXFj69d+iVi5pG6L2bRVH2qH+1rYPre73clIlXqx5lazVWpbdOGNWQppVdQlQeoIAZcL4Kg+YAPASyvmqchYCiqIoiqIoyh1GBZAPTx3yimazmQkhRJ1OJwkhpPP5PCWinoh0rbV9Zt4JIewVRbHDzANrbd85N/DeD6y1/U6nM9jZ2dn74Q9/uLe7u5taa20lbnAtdgBAQ/BYEyvOEzcu+v2+cBWB4m1f4K7DS2JLWDBpj7fCY9Xfw3w+z4+Pj+fT6fTk9PS0B2ACYEpEU2buG2PGzDy21p4RUY+ZT0MI46IopkQ0BTBN03SeJEnGzCZJkuxPf/oTPv/8cyflAXfX34+CtTaEEAoAWZIkMwDjJElOAMTW2m4URT1r7YSIMhFx3vs6NFn9QnvvzxflFlJ7gtQGi4aBhLhMjk6ghv2jyhUiUuYOaBjYF9eZhmGJ1hIFy6phfLn0Na8Xv9Pil2nNu56wTQPWSqnnKR0XTW2LJgtjWVtDoEaP4g1lb5y0eT7COQZrQRk4cwvrJW4wybVmWh5zq+rPRiNis5G3nMs08bzj8rJC2nq9q0nQN9a6pgdc9wZdtGD5rSXYXChAbPhhKfyszrA66yaxgzeKIOdUtdbO988GQec8z6r33a62Rf8a6yM+f39cB9uKva79uertvVLDUsheu9Zh5belYFkJm+1r+OJj/Z7SvEe3hfC1djSWD837CADUXv1VG0JTLAEQWmLs1nuMoiiKoijKHUIFkA8LHR4e8pMnT/jXv/41j8fjiIhSEemOx+Oe977HzIMoinaSJNnpdrv71tp9EdnN87znnOsWRdHz3neNMb3d3d3+/v7+TkUSRZE5L0TVtmlbG6sPu2t80N53l+A80aEtjlhrnYjMh8OhzbIsttZ2rbVzY8wsiqKZtXbKzBMAZ0VRnM5msxPv/amInAE4c86NjTFTAFMRmWVZRiEE/OlPfwIAuesJ0p8+fSovXrzw//Ef/+E7nU5ORDNmjgEkzrnYGNNj5n4IYTyfzydnZ2czZk7TNEUcx8YYw3WoOEX54LTFj2bv3dojpD2O6jq/kui6+r15/Zeqh2j9ZWGtbhR0kYvAW67T+1x+q0fGFevY7tlx+dK3Lr+pjLUwUXz1Tb92LyOA1+9xBAB8ceHniiAb41etHl+Lw+eibXbLn0veSQC5yMhYn9Nr81xUa7P7+fvafuvnv9TVyfqcW2kJq9QyCi9qumgbVMKLYH357WXcBOe04QafN9/6urKNC/bHtfJe9+sWpbZR77qg3Rhvq9jnXPdWRelaLGnNu3Y9WG7f5qnUPN5rqYOoDHNFVAoezfu/VHl2FsLHrThXlDa37Z1UURRFUW47KoB8OOjw8JC/+OILjuPYjMdjO5vNEmNMZzabDZh5x3u/473fS9N0v9vt7j9+/PgHvV7vsbV21zmX5Hmeeu8T730CIO12u+n+/n631+t14jiOjDHmpldSub10Oh3jvef9/X0yxtjhcNg1xuTGmNxamxtjMmPMLM/zycnJyYn3/s1sNjt2zp0Q0QkznxhjTouiiAFYYwx1Oh3p9Xr49a9/LXWC9C+//FJQhg6+UxARnj17JkmSuBBC0e/350RkiqKwImJFpAugn+f5yffff38KYGc+n8d7e3vY3d1N0zQl3Ik+ysp9ZsXIQcuepYTaqFHS9BjZUMjG6WvT2j1g3xfvy/jytnH+mzSMRu/UlLUJV1nn6xCfqjK2GOLeurxLz4sLLONYFfXuK9vWr7nu291kbogL9slVwhTVM21cpyvs+w3CS7tN9/xIugauUdS+aH88JFreHpffwhfdlRsbub3rqDVv8zmh2VFicT+TlfkURVEURVHuAyqAfBhWxI9er2eLoogApFWooZ2iKPZFZCgiHxljHnc6nR/u7+//eDgc/rDb7e6GEIz33tY5PkTEWmtNkiRRkiSW6B1jhSj3HmMM93o9y8yd4XAYOec8M/s6cToReRHJp9PplJmPT09PX0+n0zfe+zdE1E+SJA0hJHmeR0RkjDGSJIn33kuWZRLHsTs6OsLh4WF49uwZ3cWQWC9fvpS//vWv4e///u+LOI4RxzGKouBKCOkB6J+dne3leX58cnLSf/ToUeyc4yRJbOUFctOroCirNGONt3qLbvVc2GCEvdGT+b4bvbHB1Pi+13mTmLClzrdvyTZvoXZT1Mi24DLbojXPpUWFy899BT7wuXnZY+Wi8+cBXFNuFR9ye9/mfVtfd1sJyi9YaDlj6/B/22unNNvQzj9ym7efshH1BFEURVGUy6ECyPuFRqMRPXnyxMRxbKbTqTXGxEdHR7U3xwDAXgjhURzHj5Ik+agSPn7w0Ucf/WBnZ+fjwWDwUafTGdRJy+uE5gCISis0MTNp6B3lIpiZoigyzMydTieq83ZUQoUQkXjvPTPPsizrPHr0KGHm7ng87uZ53pnNZkkIoUNEHWbupGkaee9ja+3YWjvd3d3NptNp8cUXX7jnz5+7Z8+e+ZcvX96lsFgyGo1weHgYer2eK4pCBoOBADDMHEVRdJZl2VlRFCdZlh3P5/NBJSbFIYSOiMQ3vQLvg/rFSkT0Jesus8VQonv09vBO++LWnpuycXQ57a1S3SttHoqIdGuP83uKbu/L89621YZraP1c9i7FriR5UhRFURRFuf+oAPL+WOT7GA6H9ujoKPbex8fHx11jTNd73y+KYjeEsP//2buX5riu617ga639OOf0u/GgCEqKEjnOvQU6I6U8yEROVYaeUl8hH4PNjxHPMxGnGWYgDZJJSnZVUmRSTsp2yjQpEo8G+nUe+7HugA2F8Y1kUQ8CIP+/qlNoCiK4G8A53b3/vdbKOe8aY/a89/v7+/sHOzs7+9PpdK/f7+8URTGy1vYu+87A9cdbXxWWiUguy9IOBgOzu7srxhgnIu74+Ni1beu6ritFpLLWliEEX5Zl0XVdparLnPNGVevpdNoSUbderyMRxdlslmezGdH12GvV+/fvKxHlv/7rv6bRaERHR0edqjbMXBPRWlVXbdsuU0rLtm0HMcaBqia6HvfvG3kx+EAIAgDfmTdl4x4A4LuC6yYAAADAS0MA8j3ZVn7IdDq1RORjjBUzV8w8qut6lHOexBinOefdnPOuqu5572/s7e3d2tvb2x2Px+OiKCpjjLvs+wJvDmZm55wdj8eVtVa89zbG6I6Pj11d176u68o51zPG9L33PWbuOefOiagionMicqvValOWpezs7LTL5VJPT0+Jns8EuS475/n+/fty586dfHR0xF3XRWYO1trGe79h5nXOeeWcWzrnRs65hpnzdWz5BQAAAAAAAAAA8DpDAPI9UFX+5JNP5OjoyK7X66Lruqpt236McRBCmOacpyGEXefcTlmWe9ba3el0uruzs7M3Ho/3hsPhuKqqgTHGMDOGCsArIyJkrRURccwsKSWq65qm0ykTke26rrTWDqy1AyKqcs4VEVUxxiLnbFXVee9NURTSti33+30aDodhNpvF2Wx2nQaj68OHD+nw8DDlnFPXdTHn3IlIw8wbZl4bY1bW2o0xphOR17oCBAAAAAAAAAAA4DpCAPLd4/v378tgMDDz+dwTUdU0zSDnPEopjVNKeznnvRjjflEUu/1+/8bu7u7O/v7+dG9vbzocDqdVVfW89+Vl3xF4I13MlBERkZQStW3LBwcHZjAY+JTSwFrbqOq4bdvher3u13Xd27bGstZaT0SmrmtTVRXduHFDnz17RoeHh5mej2+8LiGBzmYzVVW+d+9eunHjRqiqql2tVo2IbJh5xcwra+1mWwGSUAECAAAAAAAAL9rOcAUAgEuEAOS7w0TPW1/N53MhIpdzLnLOfSIaMfOEiHaIaC/GuJ9SestauzeZTG68++67u/v7+6PpdDoYDAaVtRY/F7h0zMzeezOdTgvnnIQQClWNIhLbth0uFove48ePfdM0vus665xjEZEQAhdFwW3b5q7r8nA4zEQUP/744/TRRx9dp1ZYxMz6t3/7t8laG+u6DlVVNXVdb4wx6+2xYeaLCpA3AjNjIDoAAAAAAMBXUFVG+AEAcDVgo/07MpvN+PDwkOfzuUynU7tYLHxKqWLmQc553HXdjqruGWNu9Pv9fRHZ393d3dvf39/d29ub7uzs9AeDQeWcM/JVU6oBXhFmJmutVFVlrbWGiJyqKjPnuq6diJjNZsM5Z2FmyTkrEXHOmdu2paIoknMuMXO01oa33347bv8+0TUKQZ48eaLvv/9+FpHQdV1njGlUtVbVTUpp3bbtZrVaNaraVVVlrLXb7nWYUgkAAAAAAABEKSU2Bh3OAQAuAwKQ7wYfHh4yEZnpdGq6rnMppYKZeymloaqOVXUnpbRXluV+VVU3+v3+/t7e3s7e3t50MpkMB4NBWVWVv+w7AvACNsawMUa890RE7uIT1lqTUpLJZMKqKiIim80mt21LKSVl5qyqXc65I6K23++34/G4++STT1RV03XKBg4PD3W9XqeiKKKqdjHG1hhTq+qmaZrNfD7fGGM2o9GoHg6HZjgc+qIojDHm+txJAAAAAAAA+F7knPHaEADgEqHS4Dtw584d2ba9Ml3XOe994ZyrUkrDtm132rbdV9UbKaWb3vuD3d3dm3/6p3/61g9+8IPdt99+ezgYDIrtO+wBrgVjjB0MBtWtW7cm77777v4777xzMBqNbjrnbsYY31LVvZTSNMY4FpEeERWbzcbeuHFDiEhms9m1ufY8fPhQ33rrLVXVFEKIKaUuxtg2TVM/e/Zs/Z//+Z+Lf/mXf5n/+7//+9njx4/X6/U6pJSu08B3AAAAAAAAAACA1xIqQL4lVeWf/exnsl6vLRH5nHPhnKu6rhu0bTvKOU+Yecd7v1eW5f7u7u7u/v7+zv7+/ng6nfYHg0HpnMO7xeFaEREpisJZa8UYQyJCTdMEVc1ElIgoEFFNRA0RrWOM9ZMnT9qiKPi//uu/wocffphmsxnNZrNrERSsVit1zmVrbYwxdsaYtuu6Zr1e14vFYm2MWcUY171er9rf3y9zzu4Pf1UAAAAAAAB43V28ZsYcRQCAy4EA5Nvh+/fvy5MnT8zOzo7LORcppSqlNGiaZtS27ZiIpkVR7PR6vd1+v7+3+9x4Op0ORqNRUZYl2l7BtSNb1lpHRKyqvF6vU845M3Nu27YNIay6rlunlFYxxk1VVW1RFEREVNf1xZdSugbzQObzuVprs3Muqmpo27YLIbSbzabebDYbIloXRVHfuHGjSyklxTNbAAAAAAAAAACAS4cA5FuYzWa8bX1lu67z6/W6VxTFsGmaSUppt23bPRHZGQwGO7u7uzu3bt3a2d3dHU8mk36v13MGE7DgNWCMMWVZFvv7+6OqqvJwOMwnJyf16enpKoSwZuaNc66JMYa2bTmlxFVV0Y9//GNS1czMVzosuHv3rn7yySe6Wq3S6elpCiFEZu5EpDXGtNbalog651yw1kYRuRZVLQAAAAAAAAAAAK+7a9OH/yo6PDzkJ0+emKIoXEqpzDkPLsIPEbmxHXb+1mQy2d/f3989ODiYvvXWW8PJZNIrisKh7RW8DkREvPd+NBoNdnZ2xuPxeKcsyx1mnrZtu5NznsYYd4ho3HXdgJlLa61LKZlPPvlEVPVKnwfMTEdHR3p8fJyrqopEFIwxnXOusdbWzrnaOdc451rnXDDGXPlQBwAAAAAAAAAA4E2ACpBvjv/hH/5BfvjDHxoicjHGMqXUzzmPmXm3KIq9sixvDAaD/b29vb2dnZ3pdDodjkajyjmHtlfw2nihHZZl5tS2bTDGDHPO45zzKsa4yTm3KaVGVZOqxtVqFZ1zqa7rRESZrkEbrH6/n4koWWtjzrl7sQpERBrvfWuMiQg/AAAAAAAAAAAArgZUgHxDs9mMf/SjH0lKyeacfc65zDn3u66bMPNuVVU3Dg4Obv7whz88+JM/+ZP9GzdujKuq8iKC7zm8tnLOknO2McYqhDDsum6SUpqmlKYxxknOeZBSqpi5aJrmiyqQ2Wx2lc8LvXPnTt7f389ElMbjcVDVwMwdM7fW2sZ7XzvnWu99JyIJIQgAAAAAAAAAAMDlu8qbjlfWtmWPFEVhrLWOmYuUUhVjHOScRznnqXNubzKZ7N28eXPvxo0b08lkMvDeIwCB150QkWXmyhgz9N5PRGSHmXdCCNOu60YhhB4zF0VRuJyzqevaHB4e8lVuhXXRBmswGOT5fJ66rosi0olIa62tjTG1iNSq2sYYuxBCjDGmnHPGQHQAAAAAAAAAAIDLgRZYL4/v378vh4eH0nWd3Ww2LsZY5pz7qjpMKU1SSjsiMi2KYjoYDCbD4XDovffMV3Z/F+A7wcxijHFVVfXG4/E455yZOTFzjDE2zLzJOa9jjDUzd0VRtCmltL+/ny577X/Iw4cP9eDgIC8Wiy/mgBhjWiKqrbVrVV01TbM6Pz9fM3MVY5Rer2ettYaZzWWvHwAAAAAAAAAA4E2DaoSXpKr08OFDJiKTUnJEVKhqycxVSqmfUhrEGIdd1w1ijKWqWiISfp5+XBwAryVjDFdV5fb29nrvvPPO6I/+6I+m0+l0x1q7e1EBEmPsE1G1rZzyF1Ug9+/fv8rXI53NZjqdTrMxJocQUs45WGtbY0wjIuuu6xYnJydnv/nNb04ePXp0dnx8vFqv1yHGmC978QAAAAAAAAAAAG8iVIC8pHv37vHh4aEURWHbtvXW2lJVe6raN8YMvPdDa+1QRPrbYEQIoQe8IYwxUhSF3dnZKYuioKqq5Pj4OKaUQoxxmVI6I6J5SmlJRHVZlpvhcGjPzs7S/v5+UlW+wvMz9OHDh7qzs5N3d3dj13WBmdu2bWtVXdV1vWya5uz09LTfNE2RUrK9Xs+XZYnrLAAAAAAAwBvoKrd6BgB4U2Bj7uUJPa/+8CGEipl7zNw3xgyNMSPn3KjX6w13dnYGvV6vFBHL6H0FbwgRYWutMcaIiJCIUHg+ECMQ0TLGeBpjHIYQFsaYNREVItJNp9P4+PFjuXfvXiaiqxqA0Gw209lsplVV5dFoFJm5SynVOed113XLrusWIYSB934wHo/7KaWQcy4ve90AAAAAAADwalyEHgg/AACuBgQgL4e3sz9c13VV0zQDVR3lnCfOuelwOJzu7u5OJ88N9/b2qqqqjIjgQQ/eFCwiRETsnHO9Xo8mk8nIOZf6/f5mvV6frlark81mcx5C2Hjv681mE/r9fiSieHh4eOVngRBRnkwmyRgTiahT1ZqIlhct8LquG4YQNimlVlUTM79WLbAuZrozM2G+OwAAAAAAwP8P4QcAwNWBAORrUlW+f/++zOdzW5alE5FSRPpN04yZeWytHQ+Hw8nNmzcnN2/eHI3H436v1yvKskQAAm8kYwx77+1oNOoVRZGrqlrP5/NxCGG4Xq8HzLzKOVfe+0ZE2vF43Hrvr/q5og8ePND33nsvO+eiqnbGmLrrujUzr0RkpaobEWlEpBORRFe4ouXrQhEbAAAAAAAAAABcR1d56PCVMZvN5P79+/Lw4UPT7/dtjLFYr9f9pmlGMcZxCGGiqhNjzGgwGPTH43E1Ho+LXq/ntr2ALvsuALxyzMwiYoqicL1er+z1ej3vfV9EBqrazzn3RKRsmqao69qllMwvf/nLa7HT3u/3s/c+hxCiMaYVkdpauxaRtYhsRKQxxnQikq7wTJOv5cXwg5kRhgAAAAAAAAAAwLWBnfk/YFu2KERkDg4O7Hq99m3blm3b9rezDMYppXEIYZxzHjJz5ZzzzjljrZVt9Qd2DOFNxCLC5jkrIl5EipxzlVLqxRh7IYSKiIqu61xVVTKdTq/8uXL79m2dz+c6n89zURSxLMuuqqqamettO6zaGNMYYwIz5+segFxA8AEAAAAAAAAAANcNApCvxh999JEQkTx69Mj0+31rrfU55yqE0G/bdhRjnIQQJjHGUdd1gxBCmXM26PcI8N+28yIkxuhjjFWMsUdElYiURFQYY1xKyQwGA77q585sNtMnT57ou+++mwaDQRwMBh0zN865WkRqIrpofxW28z9eiwAEAAAAAAAAXg7eSAYAcPkwA+QrzGYzJiJDRLbf77vz8/NKVQchhFHTNBNmnlprpzs7O9PBYDDd3d0d9nq9UkQs41EO4Auqyjlnk1JyKaVCVStVrWKMlYgUqupyzlJVFd+7d4/piocGd+/ezZ999hk/efIkVVUVQgjN+fl5k1Jqcs61iLTMHF6HFlgAAAAAAAAAAADXFSpAvtxF6yspy9LlnAtm7hHRYFv5MVbVSVEUkxs3bkxv3bo1eeutt0bD4bD03hsEIAD/k6rFqt0BAAAgAElEQVRKSsnlnH1Kqcg5lznngog8EVljDB8dHV2cN1f5/FEi0g8++CAbYxIRRedcIKI259wyc8vMnYhEZs6qyD8AAAAAAADeVCJC1loqiuKylwIA8EZCBciX2FZ/yPvvv2/qunZEVBJRv23bERGNQwgT7/2k1+tNb968OT04OJjs7u6O+v2+996jAgTgBarKqio5ZxtjLFJKJREVOeci5+yIyMQYr00gy8w0m8304OAgT6fT5JwLbduGGGOnqt0L1R+vzQwQAAAAAAAAAACA6+babDhehp2dHT47OzObzcatVqsypdTPOQ+6rht1XTdMKQ2ZedDv9/vj8bg3mUyKXq9nnXMigm8twAVmJmbmnLNNKTlV9dvww+ecXQjBOuekqqrrEhzqbDbT6XSab9++nUQktW0biSimlGLXdWG9XneLxaJdLBbtZrPpQggp55wve+EAAAAAAAAAAABvCuzSf4kHDx5wjFHW67Vp29blnMsQQr/rumHbtqOu64YhhEHOue+cq6qqKqqqcs45u00/rstGLsD3bjsDRFTVbFtg+W344VXVWWtNjFG893x4eMjXpW3Uw4cP9dmzZ1lEUowxhRAiM4f1et0dHx83jx492nz++eeb4+PjpmmaEGO8HncMAAAAAAAAvhVmJlXF3hAAwCVDAPIl7ty5Q4vFgtu2NSEEV9d1Udd1r23bfgihH0LotW1bppRcjNHknPGgBvDVWFWNqlpVdarqiMjmnG3btvYiALnsRb4Enc1menR0pMfHx9l7n0Qk5ZzTfD7vHj16VP/bv/3b8j/+4z+Wjx8/3iyXyxBjTJe9aAAAAAAAAPj+qSqLCEIQAIBLhgDkSzx8+JCJSLquM0RkRcR1XVcxc7+qqsF4PB5Mp9P+cDjsee+9iBg8qAF8uYs5IERkVNUSkcs5O2a2qmqcc+Kc4/39/Wt1Ht25c0eXy6UycyaiTER5tVrF4+Pj9ne/+139+eef16enp23TNCmlhAoQAAAAAAAAAACAVwQByJd4/PgxbzabixDExhh9zrk0xvSrqhq+9dZbw4ODg8GNGzd6/X7fW2vxvQT4Ettw8ItB6NsKEMvMNudsiciklMRay0RE9+7duy4hiBKR/uVf/mVm5py2mqaJi8UiHB8ft/P5vF2v113XdSnnjAAEAAAAAADgDSIiZK297GUAALyxcAX+Cr1ej0MIQkQ2xuhTSlWv1+vv7OwM33nnnen+/v50MpmMR6NRUVWVZb4ue7YAr56qckrJ5Jy/aIOVUnI5Z2uMMSklqetahsMhHx4eMj2fo3MtAoPPPvuMTk5ONMaozrmUUkpElJg5MnMioszM1+K+AAAAAAAAAAAAvC5QtfAV6rrmuq6laRqTUrI5Z09EhbW2dM6VzrlSRHzTNGaxWPD5+TltNhuNMapelynOAK8AM5OISFEUttfrFYPBoKiqyjvn7LYFlogIExFVVcVERNflFGJmffLkiRZFoUSUt1UeeXs7q+pFayylaxLoAAAAAAAAAAAAvA5QAfIl5vM5X1SAlGV5EYC4EILvus61bWtXq5XEGEVViZmpLEudTCY0Go24qipCRQjAc8zMxhjp9Xp+MpmUzFx1XVdsW2GZnLPknL9ogXXnzp3LXvJLOTw81J///OdqjNGu614MQdL2o6ICBAAAAAAAAAAA4NVCAPIV2rbloig458xEJDlns1qtOIRAi8Wi8943IlKnlLy1lnZ2dvgHP/gB/9Ef/RF570kEBTYAREQiwmVZ2ul0Wjrn8mQyadbrdbVYLFzTNNJ1nYQQeL1e83K55GfPnvGnn356bVpg3b9/n95++20VESUi0ufythLsogIEAAAAAADgG2Pma1MpDwAAcFUgAPkKXdexMYaZWYwxknM26/VaVqsVPX36NKaU2pRSG2OUqqrMrVu3tN/v897eHk0mk8tePsCVwczsvTej0agoy1IHg0G1WCyKlJLtuu75SSbCm82G//zP/5wePXpEd+/epdlsdtlL/1pu376tZ2dn1LYtGWNURPILrfAuqj/wSgUAAAAAAF7ai8EHOk0AAAC8HAQgX8NFBQgRSdd10rYtnZ+f581mk7quiznn1O/3VURosVhQ13WUM97wDXBh2wLLGGOM916ttUVKyXnvjTFGLgIQYww/evSIf/KTn1z2kr+V56M/vqj+wEggAAAAAAD4Ri4CDwQfAAAA3wx6NH1Nqso5Z1FVUVUhoi8GNV8cL/4ZAL7a9pxioi9CxmtvW/2hRM+HoxMR5ZwvbmMOCAAAAAAAwBtEVV+L17oAANcZApA/YLPZsKp+caSUOOf8xXGxiYvgA+CbuXhC6L2/7KV8J1JK/2MWCEIPAAAAAAD4LjEzKkKugRfDj5QSfmAAAJcEAchL2D548cXH7XHxOVR/ALyEi1CR6PWoANlsNhpjVCKilBLa4AEAAAAAwHcK+w7X0+vwehcA4DpDAPLN8O/dZpQ1AnwzF08GY4yv1TnEzKj+AAAAAACA7xUqQa6P1+01LwDAdYEA5FvYvusCvf0BvqHXNTi8uB6gNB0AAAAAAAAAAODyIAD5ZvT3PmKTE+AbeJ2DQxFcXgEAAAAAAAAAAC4Tdui+phfa2bz4kYjoi4HHCEEAXt7F+ZNzfm3CEBG5uBgwEa4NAAAAAAAAAAAAl8Fe9gKuOhHRi/BDRLIxRo0x6r2nnDOJCKWUuCgKcs6RtRabnQAvSUS06zqqquqyl/KdeXHIOwAAAAAAAAAAALx6CEC+BhFREVFVzWVZ5qIoaDAYSM7Z5pxdjFHKsuSbN2/SaDSioijQ/gbgS2xn5xA9r6LKqqopJRIRWi6XNBgM6JNPPqFPP/30Mpf50nq9HuecWVVp+5FFhPi/E1GEIQAAAAAAAAAAAK8QApCv4L1XVdVtAJJVNZVlmauqotFoZIui8MaYIqVkrbWys7PDN2/epF6vhwAE4A94sa2ciKi1Vq21Wte1XudKEGMMp5R4G3zwRSUIM7+2Q98BAAAAAAAAAACuIgQgX4OIqDEm55zzaDTKu7u79N5777mdnZ2y1+tVOWdhZinLkofDIQ8GAzLGXPayAa60bSWIMrPqC2UhF+7evauz2ezVL+xbsNYyEbGIcIyRiYgvXPbaAAAAAAAAAAAA3jQIQL5CURSac84ikpg5iUgUkWitjdbaVBRFHgwGuSiKixkgfDEHBBUgAP9t2+YqxxhT27ZN0zTNer3uuq5LRJSstdkYk9u21ffee08fPHhwrQaiP3jwgH/wgx9wXddfBB7WWs45CxGJqgqqPwAAAAAAAAAAAF4tBCB/gLVWnXNZVRMzR1UNbdu25+fnjfe+EZHOe++LopCqqgjv9Ab4/6mqhhDScrns1ut1vV6vN+v1ummaJqSUsojklJL2ej198OABERFdp1Ppzp079POf/5ystayqnHO+CD0MEclFO6zLXicAAAAAAAAAAMCbBAHIl5hOp1oUhVpr88X8DyIKbdu2p6enzfn5+fr4+Hi1t7fnf/jDH/a991KWpb1Om7YAr0rOWZumiWdnZ/XR0dFysVgsu67b5JzDNly8VhUf/5uyLDnnzG3bChHJRQjywm1cHAAAAAAAAAAAAF4hBCBfYbPZ6M2bN3MIIRFRZOYuxti2bVt3Xbfpum6jqtWtW7d8jLG47PUCXFWqqjnntNlsurOzs+b8/LxOKbVFUQTvfSSiLCI5hKDvv/++fvDBB9cmEFFV/pu/+RsZDoeScxZrrVhrjTHGe+/L3d3dcjQaee+9McagNx4AAAAAAAAAAMArggDkS9y6dUuJKBNR9t7HnHNHRE0IoY4xblar1ZqI6n6/33ZdF3PO+XJXDHB1qSrlnHPXdaGu62a9Xjeq2hpjgrU2GWNyzlkHg4F+9tln9Pd///dERNchBOF79+7xrVu3uG1bzjlLCMEMh0M3Ho/L0Wg02N/f7+/v71e9Xs8iAAEAAAAAAAAAAHh1EIB8hX6/ryGEzMzROdcRUZ1S2sQYN9ba1nvfOeeCMSaJiG7b+KDNDcDvYWZlZjXGJGZOIhKJKIhIZOZorU3OuRxC0D/7sz/TJ0+eXPaSv7bDw0MeDAb8i1/8QhaLhRCRTKdT//bbb1cHBwfDyWQyGo/H/cFg4J1zCEAAAAAAAAAAAABeEWzGfYkHDx7oer1WIsplWUbvfVcURW2M2Vhr19bajbW2uQhAXocZBgDfMxWRZK2NzByYOYpIYObEzCnnrCEEJSK6e/futTifZrMZ7+/v829/+1sTQjDGGMPMtqoqN5lMiv39/d7u7m41Go3KoiisiOCaCwAAAAAA8Prj7YxYvEkWAOCSYTPuq+Wu65IxJhpjOiKqnXNra+3aObf23m+sta21NooIWmABfAURydsjbo9wcZuZUwghj0YjPTo6uhbhh6ry4eEhHx0dibXWWGsNM1tVdd571+v13HA49MPh0FdV5ay1RkTw5BcAAAAAAOD1xkTPXzNe9kIAAAAByJe6ffu2npycaFVVKeccrLWN935tjFlaa8+dcwvv/bosy41zrjPGpMteM8BVddECa9v+Kjjnum31R7DWBiJK1trcdd21CD+IiD/66COZz+fyzjvvmLIsbb/fdyLinHMu5+xyzlZVBU96AQAAAAAAAAAALgcCkK/wox/9KE8mkzQYDEKMsVPVjTFm5ZxbXhzGmFVKadM814UQLgaiX5eNXIBX5aIFVhCRYIzptrN1IjMna21++vQp3b9/n7alwlfWbDbj27dvs/feHB0d2ZSSSyl5Y0zBzF5VXUoJAQgAAAAAAAAAAMAlQgDyJe7evatPnjzRd999N202m0hEbVEUG2PMylq7LIpiaYxZENGiaZrFcrlcLZfLTdM0bUopqSoCEIAXbIegX8z96IwxrTGmE5FgrY0hhFzX9bU4b+7evUs//elPeW9vT1arlS3L0jFzwcyFqhYpJX9RAULo+QoAAAAAAAAAAHApEIB8ie1Q8/zb3/42xxgDEbW9Xm89GAyW3vvzXq93Zq2dN01z+uzZs+Pf/e53R48fPz49Pz/fdF0XEIAA/Ldt+6ssIhctsFoR6YioK8uy895Ha22eTqd6+/btq37u8L179+Sf/umf5NmzZyal5EIIhXOuIKKSiMqcc5FzdtsABAAAAAAAAAAAAC6BvewFXGV3795VIko/+9nPyHuv8/k8e+9Nr9dzTdOcE9G867rq2bNn5Wq1cl3X+aqqzHA49KrqL3v9AFeFqhIzZ2NMsNa2ItIQUWOMuQhCovc+7+/vX4QfVzYEmc1mfHBwwERkyrK0qupDCFVKqUdEPWbuqWqhqg4VIAAAAAAA8F1hZvr991rivZcAAABfDe9O/goX71p/8uRJ6vf7YX9/vxuPxw0zb5xzK2PMeYzx7Pz8/OT09PTk7OzsrG3bTc45ogIE4L9dnEtEFEWkE5HWWtt47xtjTDcYDEJRFLmua90Gj1fadDrlGKMsFgu3Xq+LlFIlIj1rbSUiFREVKSWHGSAAAAAAAPBtqOoXB9HzEORiZiK2HQAAAP4wBCBfw2w204cPHyoRpaZp4rZlz0ZVl8x8xsxzETlzzi2MMY2IxG0LLQDYeqECpLHWboioVtUm59x1XRe99+nGjRv5qp87Dx484IcPH4q11hCRU9Wibdt+jLGfUhrknHsxxirn7HPOBgEIAAAAAAB8ly4CkYsgBAAAAL4cApCvR2ezWX748KFuB5x3IrIxxixF5FxEzowxcxE5V9V1jLENIcTt/5vpCrfzAfgeqarmnHPKOYecc0fP215tmLlm5tpa25Rl2VZVFZqmycvl8qqfK3z79m0+ODiQEIJtmsa1bVuFEPoxxoGq9nPO/ZxzuR2EbggtsAAAAAAA4DuCqg8AAICXgwDkJcxms9x1XXLOhbIsa2Zeqeq5qp4x81xVT9u2nS8Wi8VyuVw1TdPEGBPaYcGbKOesKaXUdV3bNM2maZpljHGpqitr7cp7v1bVOsbYMnMYDof5stf8NcnZ2ZmJMVpmLkIIVdd1gxjjKKU03AYgX1SA5JxxnQUAAAAAgG8NWwsAAAAvDxtzL2k6neZHjx4lIup6vd6GmVfGmEWM8XyxWMw///zz40ePHj37/PPPT05PT5chhC7njGcp8MZR1ZxS6tbr9XI+n89PTk5OVqvVPISwIKL1tg1WMxwOW2ttHI1G6ejo6EqfK3fu3BEiEu+9EREXQihSSlWMcXBxqGo/pVTmnJ2qogUWAAAAAAAAAADAJbGXvYDr5uHDh/rTn/40/upXv+pSSrUxxqpqGWM8Xy6X867rjs/Pz/vr9dqpqlRV5UXEEhEzM4sIEVriwOtLt/1oNcYYm6Zpl8vl4vz8/HSxWJzEGM9UdSEiq5xzXRRFQ0TdjRs3wrNnz/J21s5V9UX7q+VyaWOMLsZYqGqVUuqr6kBEBt77nrW2FBFPRIbRmBcAAAAAAAAAAOBSoALkJd29e1d/9atf5du3b3dlWba9Xm9DROsQwqqu6/Ozs7PTo6Oj45OTk+PT09P52dnZcrlcbpqmaXPOEe2w4HWWc9YYY2rbtluv1/VyuVytVqvz9Xp9ulqtTruuO4sxLoloXZblxlrbjkajLoSQDg8P8927d6/s+TGbzfjw8FCstSbnbEXEqarftrsaGGOGg8FguLe3N5xOp/1+v18654yIIAABAAAAAAAAAAC4BKgAeUnMrNvB5vTgwYOubVvjnNvknFc55/MY44CZe8vlsjg6OnI5Z7+zs5N3dnaG0+m0X1WVWItvO7yecs6567qwWCzqxWKx2Gw2Z3Vdn7Rte8LMJ8aYuTFm4b1fiUhtrW1Wq1U4PDyMRKTMfCUDEFXle/fuyXq9FhExxhiXc/aqWnZd1xORflmWw93d3dHe3t54d3d3uLe3V1VV5YwxCJoBAAAAAOA7hUJzAACArwc78d/ARQjy8OHDVFVV8N43xpgNEa2KolgQUb9t2/L4+NgvFotivV5TSomLorDWWmOM4edfhonQDgteIznn3LZtWCwW66Ojo/PlcnkqIqfOudOiKObGmIUxZmmt3ZRlWQ+Hw05E4ieffJJ/8pOfXNkh6Pfu3eODgwPe29uTx48f25yz3VZ/FDnnkoh6ZVn2d3d3B+++++5wd3e3PxwOy7IsrbX2tTnHUcAGAAAAAAAAAADXCd6Z/A0xsx4eHibnXEwpBWtt0+v11t77hbV2HmM8XS6XJycnJydHR0fz4+Pjxenp6WaxWDSbzSbEGBOGo8PrZjv4PDRNs9lsNufL5XLetu1pzvm0KIr59vzYGGOanHNXVVU4OTlJn376ab6q1R+0DSnbtpVnz56ZGKOtqsrFGIuUUplSqkIIPWauyrIsx+NxOZlMfL/fd845ue4tsLYzXRB+AAAAAABcAaj8AAAAeDmoAPkWtgOb08HBQei6rlXVjbV2EWN0ImK7rrMppWKxWNiyLJ0xxscYuW1bmk6nRVmWF0PRAV4L2xk3UVXrnPMypTQnolNmPmXmM2ZeOuc2bdu21tpwcHCQDg4O8gcffKCz2eyyl/+lDg8PmYjk+PjYEpHruq5g5oKIyhhjKSJFzrlgZu+cs9Za45zDyQ0AAAAAAAAAAHCJsEH3Ldy9e1cPDg60qqrove+KotiIyGI75+DUGHMqIqchhNPj4+P5r3/967Nf//rXy2fPnm22VSBXtuUPwDchItkYE621tXNuaYw5Z+Y5M89F5Mx7vxSR2nvfeu/jNkS8srM/iJ5XQMzncxmPx1KWpd3O9fDOuYKISlUtY4xFjNHHGG3OGddVAAAAAAAAAACAKwAVIN8CM9PHH3+c1+t16vf7XV3XpqoqaduWY4xijDFE5GOMJsZoNpuNsdaStZbKsuSUkqaU1HtvrLUsKAeBa0hVk6qmGGNommbZdd2Zqs5F5NRae+KcOxWRubX2XFXXMcZGRML5+Xlq2zYfHh5e2fCD6Pn8j8PDQ04pGeecbZqmEJFSRHr9fr9XVVXfOTe8ceNGfzgclt57c93bXgEAAAAAAAAAALwOEIB8O/rw4UM9ODhI/X4/hBDEWktt25IxRowxTlVLVbVd19mcs10sFsZ7L957SSlpjJEmk4kvy9J67y/7/gC8tJxzjjF2m81m1TTN6Xq9Pm7b9lRV5977+bb11XlKaVUURe2ca1U1VlWVDg8Pr/Lsjy8MBgPOOZucsxMRn3MujTFVr9fr93q94WAwGO3s7Ax3d3cr771lZoSZAAAAAAAAAAAAlwwByLd09+5dvX//fn7//ffjZ599xs65bIzJzMzWWisiPqVkmNnEGE3Xdfb09FSappHVaqVN04i1Vqy14r03l31/AF6Wqsau6+rFYnF6fn5+tFqtPg8hPMs5H3vv5865M2vtwjm3cs41RBQODw8DEaXrEH4cHh7y06dPWVWtiLiUkieiwlpbTafT/s2bN0e7u7uT4XA4GgwGvV6v56y1qAABAAAAAAAAAAC4ZAhAviVmVlXN9+/fJyIKIYSsqlpVlanr2omIt9YaZjbMbHLOtmka3gYfPBqNXAjB5Zzxs4BrQ1VzzjnlnFPTNJvNZrNYrVYn6/X66Wq1eioiR0R0ug0/lsaYdVEUDRF13vtARJmIdHtcaQ8fPuQPPvhAjo+PjTHGXlSAMHNZFEU1GAx6u7u7vV6vVxVFUVhrhZkRgAAAAAAAAAAAAFwytGn5DjCzfvTRR/nJkyep3++H9XrdOec2RVEsjTFnInJqjDmy1j5l5qdd1z3bbDbHdV2fhRDWOeeLDWGAayHnnLqu69br9Wq5XM4Xi8XxarV6utlsPm+a5vMY45Ex5sQ5d+a9X/Z6vU2MsfXeh0ePHiUiysx8LX7nP/zwQ6rrWvr9vlFVp6qFiJRE1COinve+Ksuy7PV6vigKa4xBAAIAAAAAAAAAAHAFoOrgu6Oz2YyISD/++OO4Xq+5LMu6KApZrVZkjFERUSISVWVmdkVRFM65kbU2iMi12AwGIHoegLRtW8/n87P1en28Xq+ftW37VFWPiqI4ttaeWGvPrLWLnPMmhNB+8MEHgYjS3/3d3+lf/dVfXZvf91/+8pdsrWVVtSkln1IqYoyltbbMOZc5Z6eqCJMBAAAAAAAAAACuGAQg3y0lIrpz507+2c9+lvb29tq6rtl7zzFGJiIKIdhtSyxnrXUi0osxVk3TsKpmel6VY0RErLVijBERweYqXDpVTaqacs6xbdv1ZrM5W6/Xx8vl8tlms3lKRM+Y+ch7f2KtnVtrF0VRbKqqasbjcSCiRER5Nptd+bZXL+C2bSWlZL33LoRQhBCqGGMvhNDf3vaqKqqKqg8AAAAAAAAAAIArBAHI94CZdTabJSKiqqp4MpnwcrnklJI656wxRi4Go4cQiu2skNg0TRtCKIwx3nvver2eL8vSIQCBqyDnnFJKTdu2dV3X55vN5ni1Wj1dr9dP67p+VpblU2vtsYjMrbULY8xqOBxuUkrdfD6PBwcH+ToMPb+gqnz//n2Zz+dmsVi4pmkKVS1jjFXXdX0R6ccYvwhA0PUKAAAAAAAAAADgakEA8j2ZzWb68ccf58FgEJ88edIxsxhjyDlnUkqqqimEEM7Pz4Oqbqy1e8w8bdt25L0fjEajwc2bN4c7OztircXPCS5dSqnbbDbLxWJxtFqtjler1dO6rp/lnI+stcfW2mdEdGaMOVPVFTPXRNSenp7Gtm3z7du3r0v4wbPZjO/duyeHh4dCRE5EihBClVLq55yHMcZR27bDtm0HIYQypWRRAQIAAAAAAAAAAHC1YGP9+6N37tzJn3zySRKR4JzjruvIey9d1xEz5xhjWq1WOYQQcs6bGOM6hDDt9XrTtm1jVVVUFAWLCFtrZYuJCBut8H1RVdWUkqaUMhFlIsoikruuWzRNc7pcLp+uVqunq9Xqc1U9YuZja+0pM59aa5dlWS6Zua7rui3LMjx69CjduXPn2sz8mM1m/OGHH8q//uu/mqZpbM65KMuyOD8/r0Skx8xDa+2wqqpRv98fOOcqZraYAwIAAAAAAAAAAHC1IAD5Hm1bYeUPP/ww/uY3vyFVVWstl2WZc86h67q4Xq/z+fl5jDG2IYQmpdQNh8OYc879fl+cc4aZuaoqXxSFFRH8zOB7o6qUUsohhNg0Tcg5B1WN1toQQjjdbDZHq9Xq6WKx+LxpmifOuWNjzGm/35+r6sIYs04p1UVRtFVVdU+fPo1EdG1aX23bXvHR0ZFMJhObUnI556Jt24qZq5xzvyzLQb/fHw2Hw/F0Oh31er1qO9cHwSQAAAAAAAAAAMAVgs3079lsNsuz2YwODg6S955EhEUkhxCStVZTSmytJWNMFpGcUiIiyk3T5GfPnuWUUq7rOu7v7w8nk0nPGGOxzwrfF1XVEEJaLpft2dnZuuu6DRFtvPcbIjpp2/Y4pfS5tfZZURRHzrlj59xZWZYLVV0755oQQptSClVVxQcPHuRt9ce1CEDu3bvHBwcHQkTWe++IqFTVKqXUa9t2UFXVcDgcjt55553Jzs7Ozng8nozH435RFG5bnfXaU9X/8REAAAAAAAAAAOCqQgDyClyEIESkP/7xj/X4+DhVVRXats3WWg0h5BBCYuaYUorM3LVt252cnHRd18Wu64JzLnnv8zYsMcxs0A4LviOac1ZVzTHG2DRNs1wuVycnJ+d1XZ8T0blzbmGtPSai0xDCsTHm4jgdDAaLsixXqtoyczcajcLJyUl68OBB/uijj65N+EFE/ODBAyYis7OzY3POXlV7IYRBznmUcx6q6qgoitF0Oh3fvHlzPBqNBkVRlM4586YEIAAAAAAAcHXgDZIAAABfDQHIKzKbzbKq6v379/Xdd99NN27cCL/4xS9URMg5R977vA07Us45tG0bVqtVDCGoqubRaKS9Xk+dc1QURWmtLZgZbXfgW1NVzTmnGGNomqZdrVab5XK5WCwWp+v1ep5zPinL8tR7f2yMmTvn5saYeVVVp0R07r1fF0VRF0XRzefz+ISLDdcAACAASURBVM///M/pzp07+S/+4i+uS/BBRM9nfzx+/FgODg7k5OTEFUVRMHMVYxzmnEdENCKioTFmWFXVYDAY9IbDYWmM8Ze9doA/CBU7APAKfZ0rDp7CwrVwHR4/v+m59L/dN5yXAAAA8BpCAPIKMbOqaqbnVRv67Nmz7je/+Y1YaymllGKMwTnXxRhra23NzI2IdCmlZj6fNyKyCSG00+l00u/3xyJS4sUjfFuqqjHGsFwu1+fn56vVarVYrVbznPOJtfZkO+T8WEROROSMmc+Lolio6qKqqnVRFLW1tpvP5+nw8DDdv39fr8vMj99369YtfvLkiXXOeWttGWMcquo4xjhJKY1TSsOUUi/GWOScjariBIRLt/+P/0jF8fH//skXNze+6vHi9zdBLvOx5UuvHtfysgIAr5kXr0R4Hv7qfFnrzav7E/iSlX1XC774fnyb30HV//n3v8bXXPzf/0uL//N/vvm/CQAAAHAJEIC8YtuNYVVV/vTTT+N7773XMHOu6zqJSLDWtjHGtiiKNqUURSSFELqzs7MmxtiklKK1NjvnxFqbVdW+sAnL9PyLv/is9YvbL/53ZiZmZhHhC6/kGwDfO93KOV/8rn3xivEimHghoNCUUmrbdrNcLs/n8/nZcrmcd103V9VjY8yJc+7IGHPknDs1xiy890tr7VpENt77RkS6d955JxJRJiKdzWbXcpfywYMHfPv2bSEiq6q+67qKiAYppTEzT51z06IoJsaYoYgUzGzoKr/uhjfG3j/+I43+/d8vexkAAADwmlNmBCBXCGbyAQAAfD0IQC7JdgM6ffzxx0pEud/vp5RSR0RdVVXBGNM2TZNyzrHruqZt23XbtmtVbaqqCt77TlWHIuK270QXImJVle3Bqir8vOzki+P5P80kImKMkbIsrffeGGPMpX5D4DujqjmEkJqmiSmlpKqJiJSZ80UAJyJ5++ecUuo2m81mtVqdnp+fz1er1amqzr33J865U+fciTHm2Dk3F5FVjHGjqs17773XnJychF/84hfpj//4j/N1rfq4cPv2bSYiISIbYyxijD1mHnrvx0VR7Ewmk93BYLC7s7MzKcuyJyKOEIAAAAAAAAAAAABcWQhALpd+9NFH+vHHH6ezszNu25b6/T4Ph0NOKdELoUSIMTZd19V1XTdnZ2drIjqtqmpAREXO2amqzf+PvXvpbeTM7gZ+znOpe5HiTd1yt8fOxGMkaswi6GR2gR1gNgGylYF8gVm8X6KpT5DF7AzkC1jbLLPwIMvAmJUVIAgcT8Zutd1uqSVeilX1PM95FyLV7B7Jt7Gt2/9n0FUii2SR3S2Q9a9zTggmhGCW69p7b4hoFY6o9ZAkiiKTZVnU7/eTTqcTIwC5OZxzYTabNc+fP6/m83ndNE2jtXZKKc/MXinllj87pVRLRHVd17PZbHbinHseQjhm5mMiOlJKPSei50qpY6XUNEmSeRzHC2Zu/uu//ssTUdjZ2bn24ceSIiLTtq211kYhhFRE8iRJumVZ9ra2tga9Xm84HA57GxsbeZIkBoPP4UrA2X8AAAAAAAAAAOdCAHL55L333qPxeOz7/T4VRUFKKSIi0lrz8gz9OoRQichssVjMDg8Pj2ez2dMoivIQQiIiifc+DiFEImK999EyFLHLFlmrIGQVhugsy6Jer5dYa0OSJGKtlW/TBeuHnnnwXTpv3bZ5CxeFCueVOq9v2zRNM5/P58+ePZscHx/PZ7NZZYxptNYtEbVa69YYUzNzq7VeMPNCRGZN00y99xOt9URrPTHGHCulJiIytdZOQgjzuq4XSZI0h4eHrixL//DhwxsRfoiI+pd/+Rd9cnJirLW2bdtkGYAUzNyJ43hjOBz279692+v1et0kSSJrrUHrOLh0CD8AAAAAAAAAAC6EAOTyrY5ehcPDQyIi2tjYoOl0Smmaitbaa61r731FRLP5fD5r2/ZYa50TUcbMqYikyyAkFpGITqtC4hBCxMwmhGDp9M9ahxAMM+u6riMiSrvd7iLP88wYE60CBhFhZj4LHNbXX9rx5Xbf5rpvfBO+YZsf6zjzRc/7Ux3XXg8zvinwePX2VTurV+Z6SF3X9bKl1fHx8fFsOp1WWutaKVUrpZpl+LH6uVJKVVrruYjMQgjzKIqmRDSz1k6VUnNjzLxpmmpjY2OhtW7jOHZRFPlPPvkk/O3f/u21P/o6Ho/Vhx9+qOI41nmem+Pj49g5l4hI5pwrnHOl1rpM07QoyzIviiLVy3QS+QcAAAAAAAAAAMDVhQDkapDxeEzj8TgcHh7S3bt3JUmSEMexe/78eZumadU0zTyEMNVaT0QkaZomZeZEKZV67zOtdbwWgiTMHIlITEQ2hBAppTSdDnc2RKSdc1HTNNHJyUlmjEkWi4VdzQhZhhhML+YbnK2vzRKhV25feemocAjhTwazrypc1u97ThBx3pHl73W0+dXh7193+0tP9j2qU75LNYSIvBRuXBRwrLZdbbO8nyilhIjC8vrAzEFr7ReLRTOdTqu6rmfe+zkRLZYhR83MNTPXq8oPZq601pXWer4KQ0IIlTGmstZWWus6iqL66OiobZqmTdPUvfnmm+E///M/5b333gv0IsC7lkSEP/zwQ0VEJo7jaLFYxMaYlIiyuq4L733pvS/bti1FJGXmyBijmVl902MD/BQQwgEAAAAAAAAAXAwByNUh4/FYlsuwvb3tnzx54qIoarvdrp7NZotOp2OJaNa2bey9j7XWq7AjZebYe5+EEGKlVCwisXPuLAAREcPMetUSyxhjRMRMJpPIOWettYaW80GWg9PV2tD0VQByFo6EEHg1YH15AI5FhJfhxllIsgpMVgfp1rZ5qdLkom3O3pxXKku+rmLkou3Oe9yLHuvbPter26yHGK8emFy+Z+u3i4hQCGH9fi9VdKwHHmuByGo9MHNYm+3htdaubdu2aZo6hLCw1tZEVFtrK2vtQilVR1FUK6UWWuvFMvyorLWVUmoRQqidc7W1tm6apu73+22e5+7LL78Mk8nEP3z4MNCybRtd8/CDiGh3d5e3t7cVnYaD1nufKKVSEcmZuTDGlEqpgogyEYlEBLNy4EpY/nImCeGydwUAAAAAAAAA4MpCAHL1rIIQFpGwu7vr33zzTXXnzh3nvW+qqmo6nU7dNI1dziGI2rZNRCSqqioOIcREFHnvo2VbK0tElpbtr0IImoi01lp77/V8Ptd1XZtlhQh77xWdDoPm1XIVgKzQOUHI+nX0SrWIUuqsEkQptR5EfO1264nHKmB49XFeffPOCTi+MQBZPeZFj/V1Ach5Lb8u2h/v/VkAsqzeoBACyYs+WKtqD1FKrcKP9dvC8mZZhiNeKeVFJDCzWwYgbQjBMXNDRK21trHWNlrrelXNYa2trbW1UqqO43ihtV6UZblomqZRSjXW2vbzzz93RNR67/39+/f9v/7rv54FdBe+2Gtoe3ubj46OjNY6qut6FSbmaZoWWZaVxphOr9fr9Hq9IkmS2BijvunPHOAnI/L9yuIAAAAAAAAAAG4JBCBX12oouRBREJHw/vvvhyiKQrfbdaPRqJlOp43W2orIom1bG0WR9d7bEIJlZuu9N1prw8zGOae11loppZaVICqEoNq2VU3TKCLSzMzee7WqAlkJIbA6Rauqj9Nj9IrWQ49X11fBwupo8SqAWA9BVtutBxqr7VeByPptq+V6WLJuPbR4NcBYPdbZG3xBsPHqNq8+13mPcV6wsrx99RrPrmNm8d7T6rplyHEWfvDabI9VGLJCa0HIKvwgIs/Mjoi8UsotL+36OjM3xpjGWtsYY9o0TZsoipokSRpjTNvtdpuiKFoicgcHB34wGPjPPvvM7+3thfF4fGNPMT86OlJ1XZuyLCMRSY0xuda6iOO4k+d5d2Op1+uVZVkmy8Hnl73bcMsxM9Hy9wcjBAEAAAC4VdZbKYvcqPPTAAAAfhQIQK4JZpbxeOy3t7fD8fFxiKLIe+99kiQNEenZbKaJSNd1baIoUm3bajqt+tDWWqWUUiGEs3CDiNSqzZWIKK21YmY2xrD3nte2I2MMhxCUMYZO8xNm7z0rpVbBgloLOc7WV+EJEZHW+ixEMMasXtMqMCHvPa+uX1ZKvBSGrD/W+vXrQgistT5bf/V51+/zahjyqq+739c9B9H5Ycj6tquqjvXqj1XAsQo7lo8T1rYN67eHEIJSahV+BCJyROSJyBtjnDHGOec8M3sRcSEEJyJusVi4OI6dc86tbrtz544risIv7x8eP34cHj58GN56663wD//wDzf6E3Vd1yrLMkNECTNn3vtCRDppmnYHg8HG66+/3h8OhxtlWXbTNLVRFCEAgct3OhPoRfiBL74AAAAAt8rqOwm+mwAAAHwzBCDXx1lrrJ2dHXrw4EHY2tryvV6PZ7OZappGpWnKbdsq7z3nea7atlXGGHbOqRCCquuajTHMzNy2LWutWSnFWmv23qvV+vIg/1nAsbq+bVuOooiYmZ1z7JxjpRSnaUqnx9OZlVLsnOMoisg5x9ZaIiJaXbdat9bSevhhrSVr7Uu3WWvJe8/OuZe2W/Hen33aM8ac/Xze+nrAsn7f9evWnRfMvHq/9VDj1X1Zd95zOedIa/1S+LG+vqK1fvUqWWYhopQKyzZYq6U/zaZ8iOPYTafTwMy+bdtQFIXXWntjjK/rOjRNE+I4DkVR+OPjY+n1ep6W80UePny4PmfkJlIffPABL6s/4rZt07ZtixBC6b3vOud6SqkNa+1Gp9MpNzY28qIokuW/CQw/h8sjQrT2JZdFiBF+AAAAANwKfDo/87J3AwAA4NpBAHL9yN7eXtjb26PxeMwHBwe0vb3Nf/jDH3hra4sPDg54e3ub4jjmjY0Nfvr0KadpykdHRzyfz3k6nfJwOKQ4jnk2m3Gv1yNrLWdZxk3TqMViwWVZUlVVnGUZaa1XB/m5rmvOsoyWQQrVdc1KKVZKcRRFZ9sURUFN05wtkyQhIqKmaZiIqCxLatuW4zimpmlYa01Jkpytx3FMRKfBCxFR27bcti0TEa1ClNX1q/XVtqvrsyyjV29bBThEpyHM6vaLBjqsP9cqnFn9/HX3Xw991rdfD2+iKBIiImOMtG17tlyFG0SnYcjprPoXoUcIQay1IiLinAvGmLBaaq29cy6kaRqMMV5rHeq6DkopsdaG2WwWyrIMVVWFzc1NqapKtre3zwarLy90g4MPIiIej8fqyZMnuq5rE8dx3DRNxsxFXdcd59yG936jbduNEEJHa51FURTFcYzflXAlrH6pnAUfIaACBAAAAAAAAADgAjiodz0JEdHasHTZ3d3lg4MDIiLa29vjnZ0dmk6ntL+/z++88w49fvyYnz59ykREs9mMZ7MZvfXWW5SmKT99+pTv3LlDk8lEOee4qioajUZ0cnLCnU6HiIhOTk54MBgQ0YsD+51O56xF1mw2YxGhLMu4qqqXBpWvWkbR8tidMYbatuW6rqkoivXX9SeVEkopNsZQmqa0WCy4rmsmIkrT9CwoISJaXU9EVBTFSz9HUXQW2sRxfLZORC8FNK9af/xVQPPqNqvr1rddXW+tpVXIsx6mrO2XLN8DqeuaQggURZEsFguKokhCCLJ8bgkhSAhB1tdXFxEJURQF77147wMRhTRNw7Nnz6Qsy0BEcnJyIpubm2Eymch0Ol0FH0RrQ81vePBBRKR2dna43+9rrbV97bXX7HQ6Tefzed62badt2673fhWAdJ1zRdu2cQhBf/NDA/z4mPnF4HMRohAw/wMAAADgFkEVCAAAwHeHAOT6Wx+WvsJ7e3unNy4/HP3ud787O072H//xH2cBSZqmPBqNKIoiHgwGdHx8zA8ePKA//OEPbK2lk5MT+sUvfkF37tyhzz77jN988026c+cOHRwcrCoymIhoPp+fVYqsQo310IToRSsorfVZ8LG6/fj4mMuyJCKiXq93dp+Tk5Oz/RaRsyBhPZwhejmAYOaXQg0RoeFwSLPZ7CysWO1vt9ulVWDzqvl8frafTdOctwlFUfRS9cn6/lRVxUopuihgIToNcpbBBnnvKUkScc5RCIHSNJU8z2UymZCISFmWcnx8TEVRiPdelu9j+OKLL2Q+n0u/35coimQymYTDw0OZTqfy6aefym9+85uwt7dH//iP/7he5UH08t+Zm44/+OAD3t/f11prKyLxyclJ0rZt4b3veO+7WuueMaafZdmg1+ttFEVRWmsTZkYAAleCiJBifnnuBypAAAAAAAAAAAAuhADkZlo/q/9PriMiWgUkdFpBQkREu7u7TES0s7ND29vbtLe3x0REv//972lnZ4feeustIiL68MMPzx60rmsqy/KloOPhw4e0v7/Pm5ubL+3UKsw4PDwkIqJf/OIXZ7d1u92zgGXdxsYGEREdHBysV5K81M7qPK+99tqfXLdewfH2228TEdGzZ8/41eqN72o0GtHh4eGfhCDWWnr+/PlL782rVkEG0elcEGOMrF7zYDCQL774gl577TV5/PgxVVVFURTRdDqVra0tWd5HTk5O6I033pCqqs6qOqbTqezv78ujR49u8iyPb21nZ0ft7+/rra0t8+zZs7goilREitXMj7quB1mWDfM8H/Z6vdHg1EaWZam5aFAMwE9t+ftciNaCkMvcIQAAAAAAAACAqw0H9kBeCUn40aNHRES0s7Nz7qG1d99992x9FZqsrO67vb390n1WYcq63//+91/72Os+/fTTl+7/+PFjfvz48bnbfht37tw5W+7v7/9ZXWSePn164W1lWVLTNH/yfhAR7e/vv/TzeuXLct/ks88+o8ePH9NHH310dv3bb78tb7755tmfze9//3tatbTa3d2lR48enVV5LNuk3Woiwu+//76azWb66OjIlmUZM3PmnCuXba963vu+Mabf7XYHP/vZz4aDwWDQ7XY3yrKMrLWoAIErgWkZfhCRhHA6BJ0IFSAAAAAAAAAAABdAAAKvkgtmgl+4Pb2Yy0vj8fjcnqQXhSnf1qvByHpLr/P827/929c+3sOHD8/Wzwsnfgrf5nnPex2/+c1vXnovd3Z2iOhFtQ9CjxdEhPf29lQURbqua2uMiUQkDSGUIYSetXYQRdEoz/NRv98fjUajwWg02tjY2CjLskyNMVprrS77dQCcWf5+ZTodhH4WggAAAAD8yPCZAwAAAK4jBCDwQ3jpgPt3DFB+kOf8rsbj8Q+1Hz+567zvPzEmIv75z3+u9vf3tVLKxnEcz2azfDn3o5em6TBN0808z+8MBoNRv98fdrvdTlmWWZqmf15vNIAfGK8tTy+M6g8AAAD4yeBTBwAAAFxHCEAA4EYaj8f8/vvv616vZ7TWkdY6mc1muXOu07Zt33t/p9PpbA2Hw/tbW1v3e73eqNPp9IqiyDH3A64qXs7+OL2g+gMAAADgtlmdcPgTnXgIAABw7eEgHwDcRExEajabmSiKYmNM4r3PQwilMWYjSZIBM2/2er27vV7vznA4HHW73V6WZaVZ9r267BcAcBERIUWnFSDMaEcBAAAAAAAAAHARBCAAcOOMx2Pu9/u63+/btm2Tuq5z730pIt0oigZFUYySJLk7HA7v9vv9VeVHGcdxetn7DvBNePV/5tM2WAAAAAAAAAAAcC4EIABwk/B4POatrS3tnLMhhMR7XzRN0w0h9Lz3g7IsR8PhcGtzc/Nep9O52+l0Bmmaplpr/D68wHqZvWDmxKUTetGDG60PAAAAAAAAAAAuhgN+AHAT8Hg85u3tbT46OlK9Xs9UVRXXdZ23bdttmqbvnBt474dKqTt5nt/p9/t3O53OKMuyrjHGKqXQ9uprIPy4Ok5Dj4AB6AAAAAAAAAAA30Bd9g4AAPyZeDweMxGp/f193ev1DBFF8/k8cc7l3vtuCKEXQuiHEAbM3DfG9NM03ciyrEySJFsGIPh9CFffsvyDmU+DEIQgAAAAAAAAAAAXQgUIAFxrq/Cj3+/rjY0NM5vNLBEl3vuciMoQQtd73/Pe951zg7quN9q2zZ1zkYgg9PgWROSs+mO9EgQVIT89ITnNQGS1jj8DAAAAAAAAAICL4OAfAFxbIsJEpN544w2jtbZN08QhhKxpmlwpVbZtu9E0Td97P1BKDaMoGmqte8xcMLMVEbS9+o7WQw/Mn7gcq+qP1X+EQegAAAAAAAAAAOdCBQgAXEsiwru7u7rf7+sQgjXGxNPpNNNaZ977koj6dV2PRGTTWrsZx/FmmqabvV6vn2VZaYyJ0Pbq+1tVgiAEuQQvSkAI4QcAAAAAAAAAwMUQgADAdcR7e3vqV7/6lT44OIiapkkXi0VmjCm99922bXvOuYFz7k4I4c4y+Ni8e/fucDAY9Pr9fhHHcaS1RgAC19CyBdlZ+yu0wQIAAAAAAAAAOA8CEAC4bnhnZ0c9efLE5HkeOefixWKRiUhZ13VPRAYiMiCiETNvWmvvpGk66vf7g7t37/aHw2GZZVkSx7FBAALXidCLeo/T9dUQdFSBAAAAAAAAAACcBwEIAFwXTEQ8Ho9Vv9/XVVVFRJQopTIRKZ1zGyLS994PlVIjrfVmmqajNE1Ho9Fo0O/3N3q9XlmWZRrHsWVmRgcsuHaWrccUv/gZAAAAAAAAAADOhwAEAK685bBz3t3dVW+88YYJIVhrbTqZTEoiKr33q/BjJCIjZt7sdDqjwWAw2tzc3Oz3+93BYFAURZFEUYTKD7gR0AILAAAA4PbA/D0AAIDvBwEIAFxp4/FY7e3t8dHRkfrVr36lDg4O7Gw2S5g511p3mqbpeu8H3vshM49CCKMoikZpmg6Hw+Hg3r17vV6vV+R5niRJYpRS+NYA154sMw9e+z8AAAAA3GwIQQAAAL47BCAAcGWNx2P1zjvvqKqqdJqm+vDw0DRNk1hrs/l83mmapici/RDCkJmHxpjNJElGRVEM19peFd1uN42iyKhTl/2yAL4/obWCD0btBwAAAMAtIyIkgk+BAAAA3xYCEAC4ktbDj+l0aq21JoQQJUmSTafTMoTQI6KB937Ytu1Iaz2KomhzOBwOB4NBfzAYbAwGgyLP8ySKImOM0Zf9mgB+EMwvSkAAAAAAAAAAAOBCCEAA4CpiIjoLP4goev78eURESdM0pfe+G0Lot207CiFseu9HWutRmqabo9Gof//+/V6v1yuKooiXba9Q9gE3EEIQAAAAAAAAAICvgwAEAK4S3tnZUb1eT3U6HXN4eGibponbtk299ykRFW3bdpxzvbZtN5l501q7WRTFKM/z0ebm5nA0GnUHg0HZ7XYTa63RWjPyD7g51oZ/MFpgAQAAAAAAAAB8HQQgAHAVMBHRBx98oPb393Wn09F5nkdVVSXOuZSICudcwcxd59yGc67fNM2mtXYziqLRqu3VMvzIi6KI4zi2WmskH3ALIAYBAAAAAAAAADgPAhAAuExMRDQej/njjz/m/f19vbW1ZfI8N1VVJUSUiUgpIp0QwkYIYeC97zvn+s65gTFmM03Twebm5vDevXu90WhUZlkWxXFsmJkv+bUB/MhemogOAAAAAAAAAACvQAACAJeBx+Mxf/jhh+qf//mf+eDgQD948EAlSWInk4mdzWax1joLIZRE1LHW9tI0HaRpeodOB5/35vP5RhRFvU6nszEajTqDwSBbtr1SWmuM/QAAAAAAgBsN53wBAAB8MwQgAPBTUzs7O0xE+t1331XOOdPtdo3W2lZVFSulEu990rZtISJdEdmw1g6TJBltbm7ei+N4qJTqzefzXGtd5HmeD4fDotPppGmaWlR+/LCYGV+srqgXtR/48wEAAAC4DVafy/H5/HoREQ4h4A8NAOCSIAABgJ8Sf/DBB2etruq6NlVVRXEcR865RCmVtW2bOedyZi7btu157zfKstzMsuzunTt3ftbtdodxHG+0bWuJKDLGRHmeR1EUGXwR+PGsghARtFy6bEIvvvQK2mABAAAAAFwb8/kcX1oBAH5iCEAA4KfA4/GYiUg9efJE//znPzfee1tVVUxESV3XqdY6Y+bCOVe2bVtGUdTNsqxvre31er1Rv9+/0+l07nY6nX6WZWUIQRGRYmZtjFEYeP7DW4UdIoLg44oROq37QOgHAAAAAHA9tG3LcRxf9m4AANw6CEAA4MfCIkK7u7v88ccf89bWloqiSC9Fk8kk1lqnIYSMiPIQQtk0Tdd73wkhdJm5l2XZoNvtDkaj0bDf74/KshxkWdZN0zS77Bd3G4kIqkAAAAAAAAAAAODawBnTAPCDG4/HSkR4b29PbW1t6b//+783RGQnk0lUVVV6cnKSGWNyrXXJzBshhIH3fjOEcNd7/5r3/n4URa/3+/03/+Iv/uIv3njjjZ/du3fvTpZlhbUWwe0lQbUBAAAAAMBPD3P5AAAAvj8cSASAP9fZJ/HxeHxW7fHb3/5W/fKXv+TFYqHrutZt29o4jqOmaRKlVFJVVe69L0IIHefchohsENEgjuNemqa9jY2NQa/XGw4Gg0Gv1yuLosittUZrrS/xtd5Kr37ZWlWBoBrkEuFtBwAAAAAAAAD4RghAAOA8Z0e81w9w7+7unnva0fb2Nu/v7/PW1hb3+31FRDrPc/3pp5/qpmlMWZZmNpvF3vtERLKmabIQQuGc67Rt2w0hbHjve2maDtI07RdF0RsMBr3BYNDvdDobRVFkaZqiWepPbP1Ms4tCELg8cjb/HGcDAgAAAAAAAACcBwEIAKzw+nJnZ4d3dnZob2+PiIj29/fPjrI+fvyYHz58SAcHB7y8TXU6HXbO6X6/rxaLhQkh2BCCVUrZpmlirXXatm3hvS+Wy9XMj27TNBve+25RFP2NjY3e/fv3N0ajUTkYDMo8z2NjDKo+AF7BzCgEAQAAAAAAAAD4GghAAG6vl4aUP3jwgLe2tvjg4ID7/T475xQR0dHREZ+cnPBoNGIioul0yn/5l39JdV0zEak4jllElDFGzWYzPZ1OjVLKyI9I0QAAIABJREFUWmsjrXVERLH3PgkhFCJShhA6zNy11nbjON4QkU7bth3nXNntdruDwaC7tbXVGQ6HaVmWybLtFeYVXSGo/Lg60AsaAAAAAAAAAOBiCEAAbqHVgPIPP/yQ/+mf/on7/b66e/euWiwW6vXXX1fOOTUYDNSXX36prLVcFIWq65qX6zSdTpVzjo0xynuvRETNZjMtIkZEjLU2WiwWCTPHy0vqvS+9911m7kZRtJFl2UZRFD2tdemcK5qmyfv9fjEcDvN+v593Op04TVN72e8VvCAiCD8AAAAAAAAAAODaQAACcMuMx2P14YcfKiJSRKQ++eQT89d//dd6MpmYoih0XdeGiHTbtqYoCtU0jVZLzjnVNI1iZrWsEFEhBB1C0E3TaGY2Silb13XsvU+WFSCJiKQiUopIx1rbzbJsYzgc9u7du9dPkqRQSiVt20ZJksRlWcZZlllUfQAAAAAAAAAAAMCfAwEIwC0iIkxEvL+/r+I41s+fP7fGGNs0jVVKWe+91VrbpmkiZrbMbLTW2jmnjTHae6+XVR+6aRpNRFopZZRSJs9zq7W2SqnIex+FEGIiikMIsYik3vs8hFBGUdQpiqLb6/V6d+7c6eV5nltrrfdea611FEUqjmNtjEFvHwAAAAAAAAAAAPjeEIAA3BKryo+nT5+qNE2N1toQUZwkSdy2bRJFUdS27apyIw4hxM65KIRgiUiLiAkhGBExRKSZ2YQQjLXW5nke9Xq9NMuyKIqiyDkXee+tiEQhhMg5F3vvU+99ZozJu91uORwOOxsbG93lnA+9DGeImTHXAAAAAAAAAAAAAP5sCEAAboHlzA9++vSpIiKttTZpmkZN0yRa69QYk9V1nTJzqrVOiSgNIWTMnCilLBFZIoqWLa6M996IiBURG8dx3Ol00p/97GflxsZGmmVZvGyLZdaWZhmmRHQauiTdbjdNkiRSSmlmVgg9ribM/AAAAAAAAAAAgOsKAQjAzcfvvfee+vWvf63efvttRUTae2/jOI5FJBORXEQKIiqWoUceQsiZOVdKpUSUaK0jpVQUQrBt21qttVFKRcYYk2VZ2ul08sFgsNHv9/M8zxMiYhFhEVGrZQhB0+ncEa2UMlEUmSiKjFIKycc1sQqpEIpcDRhKDwAAAAAAAADw9RCAANxw4/GY33nnHb5//76az+f65OTEWmvj6XSaGWMKEemISCeEUIYQCu994b0vQgiltTZdXhKlVCwi1ntvnXOmbVvjnLNFUSS9Xi8vy7Kb53mW53m8eu71tlbLIISXB9GZmVkpxaj8AAAAAAAAAAAAgB8DAhCAm423t7d5c3NTzedzc3JyEsVxHM9ms0xrXRLRBhH1lpeOiJTe+zKEUIhIYYzJy7LMe71eniRJrLW23nsdQlDee+2911EURXmeR0VR5HEcR1pre7kvGeD2QHwIAAAAAAAAAHAxBCAAN5iI0O7uLv/d3/2d+p//+R+TZZlt2zZWSqXMnLdt2w0h9L33g2UVSEdESmYuiKiw1hZFUZTD4bAsiiK21ppVJcdaRYfWWuskSawxRl/2awa4LV6EH2iDBQAAAAAAAABwHgQgADfcO++8Q8+ePVPD4ZAnk4nWWhtmtswcaa0T7322nAFSKqVKa20niqLSWtspy7LsdDpFWZZ5nuextVYTvWhttbTezgonpAP8VJiI8E8OAAAAAAAAAOBCCEAAbrDd3V3e2trihw8fktaai6JgEeHFYqGdczqEYIkoWl5iZk6stVmSJEVZlp2yLItut5slSZJGUWS01qjwALgShIh4OQQdIQgAAAAAAAAAwHkQgADccA8fPqTXXnuN2ralZ8+eUdu2TESklFIiophZEZEWEcPMNkmSqNfrZcPhsMzzPE/TNI6iyCy3A4BLxmvL03W0wAIAAAAAAAAAOA8OaALcYI8ePZLJZCLeewkhSBzHwRgTlFJeRFpmbpm5YeaWiFZLx8xOKeWYOSwvwsw4ygpw2ZhftL16kYAAAAAAwC0jImcXAAAAuBgCEIAb7t133xXnnDjnwvPnz0Nd105E2hBCQ0QLEVkQUbW6hBCqpmnm8/l8XlVVVdd14733gk/WAFcPZoAAAAAAAFwL1lp8pwYAuARogQVw88l8Pg/OOc/MLoTQ1nXdKKUWSql5CGFCRAkRae+9Xs4HUXVdc1mWod/vizFGG2O0UshMAS7dMosUERSAAAAAANxSjBNhrhWllHjvKcsymc/nl707AAC3CgIQgBuMmUVEqKoqaZomKKWcc65l5rpt24VSasrMVmtttNYhhODbtnXOudp7vxCRKo7jeZ7nldY6FRETQmAROWu+s1oXEWZmCiEoEeG1i2JmVkopa60yxiilFDM+sQP8WZb/AAl9sAAAAAAAri60kwYAuFwIQABugU8++SQ8ePDAV1XFVVWpuq5ra60OIZhlcBG01nUIoXLOTZ1zx3VdHzPzUZIknSzLuiGExFprRUSJiFoGHWcXIlIhBL26OOfMaqmUMlEU2bIsbVEUNo5jjfwD4Pt7EX4QYQg6AAAAAAAAAMD5EIAA3HDMTOPxWI6OjuT111/39+7daw8ODpS1lubzORtjPBE1bdtW3vupUupYKZUxc+a9z6bTaa6UyqMoipVSVkR0CMGEEIz33hCRXq0752wIwTrnorZtY+995L2PlFJxp9NJ7927l1lrlbVWKaWQgAAAAAAAAAAAAMCPBgEIwM0njx49or29vfDHP/6R0jT1cRw3q76jWms3m81a7/3CWjut6zrRWicikjjnkqqqYu99YoyJmNkuQw7jvbciYkXEeO/Pgg/nXLy8pM65pG3bxFqbtm2b53nusizzWuskjmNrjNHMrNAOCwAAAAAAAAAAAH5oCEAAboHlLJCwu7srb7/9tlRVJVprUUp5Imq9940xZh5CiJZtriLvfRxCsIvFwk6n00hELBGthx5RCMGurm/bNg4hxCGEuGma1DmXhRCStm0za22mlCrLsmyTJHFKqTaEkGZZlmitLQIQgG9HBO2uAAAAAAAAAAC+LQQgALfEavDaeDwO29vb8vOf/zx8+eWXLs/zhojqLMv0dDo1TdMYrbXJ89w0TWO89zaOY+O9t0op0zSNZWazDC6Mcy4SEds0TeSci733cRRFaV3XmXMuNcZkRJTXdd356quvJs65blVV3dFo1FNKqTRNtVJKXe67A3ANMRMGoAMAAAAAAAAAXAwBCMDtIuPxWIiIx+OxPHr0yBMRv//++85aq4hIj0Yj5ZzT3nttrdWdTkeHEDSd/r4wTdMYZjZEZJjZ1HVtQwjWWns2+8M5lzBz6r1P27bNQgh5CGFycnLSaZpmTkSLKIpCnudKax2IKNFaayLSqAYBuNir/zhQEQIAAAAAAAAAcDEEIAC3k4zHYxmPx6ufvYisTifnjz76SHW7XfX06VOV57mqqkpnWaattappGt227WrwuV4sFmfBSF3XURRFtq7rmJlT51yitU6bpsmapinruu5WVTXXWtdZloWyLJmZfZ7nPoqizBjDRKQv600BuMp4fSlCqP8AAAAAAAAAAPh6CEAAgIjOWmSJiPDDhw+FiMLx8bEyxnBVVf7evXt8eHioJpOJSpJEJUminj17ppumUVEUKWOMVkrpuq6Ncy4yxkTe+1hrHRtj0hBCycwTrfXMOTd//vz5whhTLxaLeb/fH3a7XVZKqWUlCAAAAAAAAAAAAMCfBQEIALzklSAkEBF//PHH/O6779L9+/f5o48+4jRNOYoijuNYTadTJiKOooifPXumsyxTIQQTx7Exxti6riOtdRxFUVHX9YyI5s65+cnJybxt26ppmkop1cZxzMzsjTEJEbGIsIgoEeElpbVWSilWSuHEdwAAAAAAuJXQBhUAAODbQwACAOdaDU0noj/5dL1sl0VvvfUWERHv7e0xEdH+/j5vb2+r0WikmqbRSikzmUyMiETz+bz23jsiapumaeq6rqfTaUNEbRzHkue5FpFGa52FEFYttkwIQWutjTHG5HlurLWa0CYLAAAAAABuGQQfAAAA3x0CEAD4ztbCkZWzwepEJP/93/8tr7/+ujRNI1rrUNe1GGM4iiLVNA0ppQIRtd57V9d1O5lM6i+++GIWx3GPiHLvfdK2beKcS9q2TeI4TouiSO/evZuVZclokwUAAAAAAAAAAADfBAEIAPy5zipFxuMxL5fy9ttvy9OnT2U2m4U8z2U2m5G1lr33wsyOiBpmbhaLxeLo6GjeNM2JUmojhFA653LnXN62bdk0TVGWZdHv98ssy9gYw8YYZmallGJmRjssuJ1wAiAAAADArbT6CoSKEAAAgG+GAAQAfkhCRDQej0VEZG9vT/7whz+Efr8vGxsbMp1OxVrr6rpulFILY0zVtu3s+fPnJ4eHh0dE1GnbtkNEpXOuE0LYaNu2u7Gx0fXet51Oh4wxnpnzJEmMtdaiGgRuo9WXXuR/AAAAAAAAAAAXQwACAD+KZZusMB6P+e7du0JEkiRJmEwmjoic1rqJoqh2zi1CCHMimnrvp8w8cc51jTEz7/0ihLBo27aZzWbtkydPgnOurarKDwaDvCxLhQAEAAAAAABuMlR6AAAAfH8IQADgxyTLahDe3d2V7e1t75xzeZ63IYQmz/OaiBZa67n3fta2bVXX9TyEULVtO2/btlZK1UqpZrFYNF988YVv27at69pbayWKIhVFkSKi015Yp2fD45R4AAAAAAAAAAAAQAACAD++ZTWIEBGJSNjd3fVbW1t+NBq1JycnbRzHjfe+XiwWbZqm9Xw+r7XWCyJqRaRxzjUhhLqu65aZG2ZuO51OSJKElFISRZE1xqAdFgAAAAAAAAAAAJxBAAIAP6lVGCIisru7Kzs7O+GTTz7xo9HIHR4eeiJqQgh127YLZq6jKJoz8yyEMPHez5ummU2n0/nTp09rImqapqnLsuwURZErpTRmIgAAAAAAAAAAAAARkbrsHQCA22k1I+Tjjz/2W1tbbVVVzXQ6rY6OjmZN05x474+iKPqKiL6MouiJMeYgjuPPReTzuq4///LLLz///PPPDx4/fvx0Op2eNE2zCCF4EQly2iQXjXIBAAAAAAAAAABuMVSAAMClGY/HgYh4PB7LO++8I0QUrLV+Mpk4a61rmsYnSdISUcPMNTO3IYTGOdc0TdMSkWdmV5YlxXEsSimx1ibGGKuUMqgGgZvqbBAmBmICAAAAAAAAAFwIFSAAcNlkPB7L7373u0BEfjQatbPZrGHmBTPPjTFTETnRWj/XWj9TSj0loidN0xzMZrODyWTy+Ojo6PNnz54dHB8fP62qauKca4koXPLrAvhxMZGg0AkAAAAAAAAA4EKoAAGAq0DG4/FqyUQUDg8PJc9zGg6HwXsfoihyIQQXQmiIqNZaOxHx8/m8Pjg4qOfzeTWfz9u7d++StdYaYyLMRIebjJf/AQAAAAAAAADA+RCAAMBVIURE4/FYiIh2dnb8gwcPqNPpSJ7nwXu/CkBapVSzDEBa59zi5ORk0bZtzcwhz3O21nLTNJ6Z4xCC1lprY4yO41gt4agxXHNMIihyAgAAAAAAAAD4OghAAOBK2tvbC0REW1tb0rZt0Fr7sizdYrFwVVW1aZr6pml8CMG1beuIyJ+cnKijoyMjIsoY04pI5r1PrLVxURRxt9uNkiRhBCBwI/BLCwAAAIAfFT5zAAAAwHWEAAQArirZ29sLDx48kO3t7XB0dOSfP3/uNjY2XFEUrVLKWWu9c84ppRwzh6qq9BdffKGOj499CGHetm3Xe98piqK4e/duiKJIRVGE2Udwba0OPDDjIAQAAAAAAAAAwDdBAAIAV5ksW2KxiITd3V2O4zj0er1grZWTkxNWSolSipiZnHPq5OSEJpOJc84tmqaZe++bwWDgO50OO+diETFEhOEgcAMwiRDGoAMAAAAAAAAAXAABCABcB8LMREQiIrK3txc2NjaEiKhtWx9CkKZpfNu2q1khi6Zp5k3TVETk0zSltm1tCKEQkfhSXwnAD0Dk9IIqEAAAAAAAAACAiyEAAYBrhZllPB7L1taWJ6Km1+tJ0zRMRCGKohBCaEMICyKqicgxs0qSxEZRlBtjWqUUJkfDNbaKPE7rPhgJCAAAAMCtsTwp7GwJAAAA3wy98AHg2hmPx3JwcOAfPnzYHh0dtVEUVVEUzYwxJ1mWHRpjvkqS5Msoip5aa78yxjxj5kPn3PO6rqdt21beeyciCEPg2hGR0wsJ2l8BAAAAAAAAAHwNVIAAwHW0mg1CW1tblOe5FEURptOpr6rKJUniF4sFxXFsRCRRSiVt26az2SwzxigRkTiOc2NMpLVGEAzXDjPjzD8AAAAAAAAAgG+AAAQArq1Hjx4JEfm9vT2eTqdUFAWlaSrT6VRCCMo5Z0Ukmc/n+quvvqKqqvxoNKp7vV49GAzuKKVYa43fg3B9rHXAYsIMEAAAAAAAAACAr4MDfwBwbTGziAgRkScimk6n1DQNKaVIRDQzR8wcLxYLHULg6XQqIsJKKRVFUUpEWkS01lorpZiZUQ0CV5bI6cwPBB8AAABwGdB68+oQEfLeU9M0NJ1OyVpL3nuKooi01qQUvtYAAACsIAABgGttGYIEIpL3339foiiSfr8vzjllrTUhBFPXNVdVJSEEr5QyxpjIGFOGEKz33iRJEltrjTH4lQhXnBAx8UvDzxlxCAAAAMCtIiLUti1Np1P66quvyHtPnU5nVRGPAAQAAGANjvYBwLXHzEJEtLOzE/7f//t/UlWVKKW40+moqqrOPv0756RpmuTZs2dJ27bFycmJHg6HajgcdpRSbIzRl/cqAL47IcIodAAAAIBbJoRAVVXRYrGgw8ND6na7dOfOHbp//z5prclae9m7CAAAcGUgAAGAm0L29vbC3t4effDBB9Lv94mIKM9zev78ubRtS9basFgs4qZpkuPj43w+n2vvvYmiSC0HSrMxRqEdFlxJTGe9J5at3wAAAADgFgohkHOOqqqiqqpoMpkQEVGv16M8zy957wAAAK4WBCAAcJMIEdF7773nP/jgA/qbv/kb+vTTTzlJEk6SRDVNw1VVZW3bZm3bFt772BiT5nluiUiFEFSe59acuuSXAnAOXlsyWl8BAAAA3Cark2BWLbBmsxk9f/6cRIQ6nQ41TUMhhEveSwAAgKsFR/gA4Eba39+Xo6Oj8Nprr7XT6bQxxlRVVRlmnlhrnxNR6ZxLjo+PIyLi+Xzue72ev3PnTlkUBdphwZUmcnpB9ysAAACA24eZzy5EqA4GAAD4OmjxAgA30ng8ll6vF7TW3jnXMPMijuN5FEUTZj42xhx67786OTn56vPPP//qs88+O/ryyy8nVVXV3nt/2fsPcC55kXmInE7/wPddAAAAAEAIAgAAcD4EIABwU8l7770XptOpU0q1VVXVTdNURDRl5uM4jr8SkacnJydPnz59+tWzZ88Oj4+PT+q6bkIICEDg6lmFH/JK4Qc6YQEAAAAAAAAAnAsBCADcZLKzsxOapvEnJycujuNGKVUlSbJqg3WotX62XB4bY2bGmIaZ0Tj3HCKCM8suGdNa72cmhB8AAAAAAAAAAF8DAQgA3GjMLP/+7/8e4jh2nU6nMcZUzDzVWj+PouiImQ+11kfW2mNjzISIFiGE1nvvQwhBcMQfrgpeVn6sDT/HX04AAAD4qeC8C4Bvh5nxMR0A4ApBAAIAN94HH3wQfvnLX/rZbOaMMTURzYlowszPrbXPjTFHSqnnIYTjqqqOZ7PZdD6fz9u2bUQE7bDgypBl5HE2/5xRBgIAAAAAcJUsz6ETZpYQ0FwAAOCyIQABgBuPmel3v/tdaJrGN03TRFFUZVk2YeYTInpujHnetu3hdDr96smTJ18+efLk6dOnTw9ns9m8bVsEIHBlMPNZ3nG6zsg/AAAAAACuIBEhpRSqQQAALhkCEAC4DWQ8HsvBwYEnovbo6Kj+6quvKmaeGmNOrLXHTdM8Pzo6Ovy///u/p3/84x+ffv7554fHx8ezuq7bcEqW7bBu1QdYZhxdv0pOTyY7DT5kFYAAAAAA/ARu1YdgAAAAuDHMZe8A/Oi+7dGxc7cbj8d/1pN/j/vjc/W3h/fqu5HxeEw7Ozvh17/+tYuiSGaz2UJrPdNaT5qmOXbOZbPZrHDORd77KEmSmJkT772NokhHUaSstTjiDJdCiEgpJhEhVkwUZDkIHX8lAQAAAAAAAADOgwDk+uNXli+FDh9//PFLR8Z2dnZof3//T46WPX78+NwjaFtbW3/Wzv3mN7/5Ttu/9tpr3+ug/vb29jfeb29v7/s89JX14MGDC1/zOcGTvLK8rWRvby8Qnb5/r7/+ehNCWHjvZ0R04pxLmqbJlFKxiMRKqbRpmmQ2m9nBYBCVZRkZYzSqIuAyMJ2W0TO9mAGCv4sAAAAAAAAAABdDAHI98XKoFu3u7vL29jYT0UvBxtbWFi+XdHBwwEREz5494ydPnlC/36fDw0N+4403zh6w0+mcexRtNpvR/fv3v9dOfvbZZ/RXf/VX33r7Xq/3vQ7OTyYTefLkyTdud/fu3e/z8ERENBgMrlRwsLW1deH+fPTRRzQej89u//jjj4WIeBmYMBHRo0ePlvOTmej2hSKyt7cX9vb2eDwe+zzPm7Is59baiVIqcs5li8UiaZommUwmxeHhYT4cDmMiojiOdZZl+rJfANxOq3+oQYQU0WkLLKVQAQIAAAAAAAAAcAEEINcDj8dj/vjjj/nBgwe8tbXFv/3tb1VZlry1taX29/dVmqbc7/d5Pp9zHMd8eHjIdV1zFEVMRFzXNW9tbdHh4SHneU7WWj4+PiYioqZpXjp61rbt2c/GGP7f//3f773jVVWde7219k8OuldV9SfXR1H0rQ7Ot237jdsNBoM/ue6ix59MJi/9XNc1ERHFcSzrt33b/fshxHF89lz/n707220kSe8F/n0RkRuTm6illq7pnq5ZbEhtwIAB35wD9DyAb+sV5jWa9Qo2YMDnEbpewgYM382FMS5dGHB7gJnp7unqKknccouI71yISSUpaquuKomq/w+QRJG5RCbJZDL+GRHffffd0n1xHC8ee/z4McVxLHmeS5Ik8vnnn9Pu7q6fTqfS7XZlNBrJP/3TP0kURX44HMrLly/lxYsX9QXlH0sYIkREg8HARVFUxHE8y7IssNYGRJRYayPnXDIejzvOubZSKnn06JGx1oYigqvu4VYsXnuN118dhgMAAAAAAAAAwHkIQO4+Hg6HTETq4OBAffbZZ0prrdM01aPRSGutdb/f10mSKO+9iuNYi4gyxrDWWjnnOAxDpbVmImKtNXvvKYoizvOciYicc4u/YRgSNbrTstY2778xpdS5+7TW52rsnHMy/7s0TVVVa6c3xizdd9F0K+tdO826+1qt1tplFEVBnU5nMf1V61ydt2l1G66zzHo/1ay1QkSU57nU4VEcx2KtlSRJhIh8r9cTInLtdtvP//dE5JMkcd1u1x8cHLiDgwP/8uVLOTg4kEbrkftesypv3rxxT58+tVmWFVrrTEQmSqnEe98qy7JdluUoDMNJWZYzEUmIyDHzoiUNwId2OuQHk3hPfn4bLUAAAAAAAAAAANZDAHK3LcKPwWCgi6IwZVmaOI5NVVWBiARKKdNqtQJm1mVZGhHRSimttdYioohIW2tVEASslGJmZu+9IiJmZvLeMxGx95611uycI+89G3P60pjfT8450vrmPf9cNI9SalG5bq09V+nffLxZ6V/f75wTa+3S9N77xe3mY41piJmXHtNaSx26rJZ7dRlKKYnjeHG/Ukquuvq6uR3rWos0H695789tb80Ys/Q4M4v3Xub7SE6fdhFjjA+CwBOR11o7770zxrhWq2WNMbYsSzsajVyaptY5Z6MosvMusvyzZ8+aLULuO398fGwHg0E5nU7zIAgCa+1EKTVWSo201uMgCKZBEMy01l2llL/tAsPHi/l0AHSZd4FFROTp43ijAgAAAAAAAAC8DQQgdw8TEdXBx+vXr/X29rYmIpMkSUBEYVVVobU2tNZGIhJ670MiCkTEMLOpqsqIiLHWGiJSIqJFhMuyVHzad48SERYRds4tbs8r1piZuaoqEhFutuCoA4ZVSqmly4+dczS/Sv5Cqy0Z6nm898TMS6GEnBZK6tvN6evpmknEPBBYV06ZBzyL8jXDjNXyrPLeL0IWZhYRWTtdc33N6VeXu+7x1fucc6thEDX3hYjIfLtkvg88EXkR8UVReK21IyLLzJaIqizLrIhUrVarVEpV1tpyb2+vyvPc7u7uuqIo3MOHD/1vf/tbf3R0xPe9RchXX30l/+///T8fhmGV53lhrTXOuZn3fqqUmiilxsw8JqJJURTTyWTSiqIoDILA6FPM6A8LPiR0fwUAAADw0cNXEAAAgOtDAHJ3sIjQ8+fPmYgUEamTkxP95MkT0+l0jIhExpiwqqrYORdba2MRicuyjEUkng/eHHrvA+99ICKBc84wsxYR7b1X85YfiojOBSHzx4nniIjqx64qeN2FVm3eT/1qzZysTrPY8Ma0zbCj/r85Tf3/6v3NYKAZcNSPra5HKSUXBSjNeVbL2Fz26npWNde7GnTM5z93/+q0zRBkNfyo/yqlvIiI1tqLiCcir5Ry3nvnvbfMbI0xZVVVpYhUYRiW0+m0CIKgCIIgH4/HZVVVZavVqsqytE+ePHFZlrkvvvjCRVHkv/76a394eCjD4XDxtFy0zZuGmWU4HDoiImtt6ZzTSqkZM0+UUmNjzIiITsqy7BwfH7eMMZFzznS73ThN00gppRGAwG2YHzCIEIIAAADAh4LzjjuhbhUMAAAA14MA5G7g4XDIL1684H/4h39Qv//97/WPP/6o4zg2SZKEeZ6HcRxH0+k0CYIgKcuy5b1vEVFCRIlzrjUPRELvfei9D51zoYgERKS990Ypxd57TY0WIfPbTKetThSfNmuo63N7u+EOAAAgAElEQVTr+4nm3WVdpNlSZF1F/7r/V6er6/PrRTZuL4Ud9XTr5muuoxkkrJvuohBjJaA4d9+61ikX7ZfLynNR6NMMOFbDjma569Yf8y69RCnlq6qqww+vlLJaa+ucs8xcEVHOzKVSqrDWFsycO+cy732otc7DMCyIqGy1WlWr1ar29vbsbDazW1tbjogc3eOusYbDoTx79swfHBxYIqpEpAjDMNNaT5VSE+fcaDKZnPzxj3+MR6ORmUwm+pNPPhFjjA7D8PwgNwAfgBdZjAfy4//9vzT+q78iNQ9E6helEiGupxMhFiKm+v+Vg3z9U4cqzNcc6KY+HFwydXPUnPnts6mZLj6kcGMKWbpH5tuxut7T+1fLsjLtYpXN9a4vf7MEqy4aDIibjy22+9yGnz0otLI9Z/u03vbz6+HF8uuPt+X1NVfRnHv9fjt9zs/fv/K0vYWzOZvlfZtlXXceXlNqaTx/61/Zq8/vu8q1r/q45JXXyM3LcGcjeHmfJws3WfJlO+i6y7nOa+Zq15lj9fW5/shzNvW5+5kXN2V17vOHxqsKs3aadSU4N9m6O675Ym0enq+a5dy0K9tef39Z/Ri6auObb8e6DPUybvTMy8XP2EWl4OYKzz2L50sgK7dlXlIhIREiaSxO5uOGLd2e/+953oycmDwJCTP5ebebVHfBSUTjv/7r628/AAAAwB2BAOR2LY3xcXR0pP/zP/9Ti0gQBEHQarVCa21MRHGe5wkRJVmWpc65lIjSKIpacRynSZKkzJwQUSgioXMudM4FImK890ZENM1bfoiImo8Norz3qu7yauUv1bcXBb0kAWmEJosrUVYCj/Nfg9ZMtyboaM67tmVIPf1Fj62btvl3JXhZvf/CMl70/6or9sNiXavbQI0QqH6sGdY0ApL5dxj2dWsQZnbzrq+cMaZSSlVa68J7XzjnijzPsyzLZlmWZcw801pnRJQZYwqlVElERVVVZRAE5dHRUUVE1dOnTy0RuYODg9PvRkR+3jXWfQhD5MWLF36+bZaZS2bOvfeZUmpMpy1AWkdHR2FRFIHWOhoMBqFzLp4HSLddfvgI1UGFiNCP/+f/ENHpQZ6ZadHUbx6AnCbfZ/cppkUYoohJzcOO06Z/p5U9ddU70yIPuV6Z5paOoc0qn5UapLO8fXm+RZV5MzPg5uOrBZpPKMsrWGxX4+G127J0JONF2WS+PD4/0Tl1mZnPpj0Lb5olbl61eUnwshRCyUowxcTzCq7Th2W+jcvh0FlZeLFb1oVPzfmWsppFMRdJy/zf80HJ2ec6rUwniyLWEy8muWCXLm/5PLRbeR2tfR7r1+4Fgc5q5eFZua/zAl9788KJLz09WFrA+tfC2pfpuvrsDx6AXPNjX5b+rLXu1PJaS7/hmcfZelZeizdexsqM0qycvrzG/vQ9djZfYw5afQ0sHUvPLUmW35eLe8+WeXbEuvgUVBbF5cb+OP8eXgoCmtuwWn654P1er2PN1i79LyvTrr7WG0EGLY41q9OelUNopTzN381lr31e1z03tAgBzta9jjT2k5wta2V/nD07F7xeVl8Di29DSwfx04BjfkA8DShOj5gyX76ns8c9MQkTCavTcIOI/DwA8cx0esWTkCUhK6c/dQAiRIsxyO5u6goAAABwMQQgt4eHwyE/evRIh2Go626r5l1YRcaY2DmXWGtT733Le9+qqipl5tRamyql2lEUtdM0bW9vb3eiKEqYORQR45wLvPfGOWfmrT1Www+ehx/1hcL1wOh1F1hLoQY1659WTnov6iLrshYgq2OJrAQeRMvfRGT1vqtaf9C5bzKXhxjN9a+WezUguaLcF65ztQXIusfXPLa0bastReZfRGQekHhmlvkg3b4OQpjZGWMqZq5EJM+yLH/16tU0y7JJlmUzrfVMaz1TSmVElCmlcqVUrrXOlFKZ1rooiqLIsqx49OhRlSSJdc65sizd119/7Z89e+ZXy76h5OXLl+7Jkydud3e3cs4VURTNiGhsrT221sZZloVVVUWdTicty7ItIpbuRwAEm6q+ivM0RCVHRKpxZacXIT3///RDgOatQ06DkTr4UKxOB1afV3JzIxBpVjZdURS6sCZ2UcF8VjG9qNBuhBqrVfP1DV6+0Vhms7K+WcF2Ft40l8VLlVdni6nDBrqgHOcDjHMbuPhTL3fxd838K59A50OH+QJk0cpnJbiRZhnPylwHNnWAVd+mxjLrNdYV/0v7Yc3tRUWq0GL5zfubu+ts+2Rp+xeVho1lnmvVslLJWi9nUe5GMLaIgJovkvnymy2Amr+lsYPP9twFrWEus7Ktl014ra5JmM6VYTk8pMb9l83/oV3vo+/iM6gz584rrzHNDYqwtlRvM+v6AOR8yHDRNjcrzJfevdcozGK+1TIstfZorH9RtrNH1pV/ddp6mtVpV197Z9M2H5/P19ioc5smy9ty0aavXIS08thKQLMalsw/w87Ws7KtJBd+pNWbve7hOlA4C1ia+3VlnqUnltfc17x1dQBST7+4R1Zew/PdXgcV9bHQN14biy8VSs0DktPww5MQsSJHctrcm4icELnGOpoBCMIPAAAA2FQIQG4HExF/++23+tGjR8Hx8XHYbrejoijiIAiSuoWH975rre2JSNtam1pr2/Of1BiTdjqdTq/X6/7sZz/rdrvdJAxDIyLKe78Y86MOPORsPA8mOg0uGuFFs+ur1XIu3/EOTnxXKwUuCxKaFf4XDcJ+nQr4lQDkwnkvCEAu89Zfwa+z7qumITptGbPaTVYdoDCz11o7ZvZ5nhfHx8dZnuejo6Ojk6IopmEYZiKSGWNm1tqpMWZGRFPn3LSqqrFzbsrMs1arNfXeZ9bast1ul1prS0TVixcvaDgcynA4XP/kbJCDgwN5/fp13X1YEYbhVEROjDFRWZbGORcEQRCHYdgJw7CvlHL3JPyBTde42nVRATKvPPciixYhiw8AorOwg4hI3KJSh5mIpVFrQrSoiF+/bmpMe36qs8rd+TWp0rxfVmt1aFGZvW5JS/M2K+Pnv3n5vtXgYTUmX25BsRp70PLEF+yBpX3DTCy0qOxvVrTTUklWt2xeWS6Nz9jVsjKR+MVqqFnBvlRuOau9qyvzFlcj1xWD8wVxcz0rm1gHJKt75aIWOOe2rLE/xdczr4Yr5/dDPbM0Xijil0vB84XXz+dyK53zZZ1v+tk+WSr06jXtV3zuX/sU6Ir9s1jZWTnWrf/cK3Fdxfp1i/ROXe+j76oK/rol21VLPvfeeetP3rf/yF57PUzj36Wr+tfWoJ+10eDlGnxaDm8vOdeeX+F/fr2rQUy93EZhLihY/dlR15Cv5iRy7sb5f89t10oLl4sCrLXPxqK4zUCl8bDQ+e2X5eBnubXachnXkpV/LmmZdJblytkd5xYhi7LJ0v5v3qgPhNcpUz1HI6FpBkgijUP/2W+Rs/CC1elFEezptBVI/TgRCXvyMm/ePf8c9SLkvT8LTxB+AAAAwIZDAPJhLbq8IiKVpmmgtY7iOE5ms1krCILEWtv23necc92qqvoisqW17gZB0FFKtYmoba1NtNatra2tdr/f7/T7/W63243DMKzH9liEG6tBR12Q1ZYbF7XkWBT8HZ/0XuvKSLp5uPFT1v2hK7OvWt+6oOiq5TRbx6wEITKbzSrvfdbr9Ua9Xq/nnJsaY4p5a49pVVVT7/3Eez92zo2VUqn3fqy1HhdFESmlJnme5yKSW2vLqqpUp9Ox+/v77uuvv3b3oTXIF1984UejkWXm0hiTB0EwyfM8DoIgrKqqpbVui8ikqqpZnud5EARJFEWstVZKKV6XIgJ8MHLaZzeJUF3nTESLKz0X44Ewk1uEH82YQJbqYnjlxtUv7ouCAqmLd1bp3qz/80vpw3Jl55rat3WV7fO0Z6nw5wOCpYepWUu/7nNhpep/zVKaYQwtKtLlrCZquZXChcuoK/wvmWYeHjQr/tcFNUutJxb1Vc37fWObV5bQ3H0rdXTNYOXcxGtKwo3fi/1Rt2q5tBL/oorfuhinr+ylbrbWlGfxil5z6fpZS5qznbkaqv0055/HS0NEaZbg4iWeS6jOLeP6mq153s76ec9VeF+1inWVx9df3Vu6+cIWIcFl889f49dac7MWf+mttVpZfurcupsBxUXFOT0bvLrcdQglSzNeaW0AQs3nvRnrXBAgX7ng81MsPReLsOOS15HQhY+vC1hOy3vZYuTCcq2WmS+4fzFHY/3XOnmcb+uiGCtlPreGOuBoTCx+/hmwaJl3+tc3N49OW+svWn4QIfwAAACAjYcA5MPhZ8+eqZcvX+onT57oX/7ylzrLsrgoisR7nzrn2t77tve+S0Rda23fe7+llBoYY/qdTqebJElHKdV2zkVKqbjX67V6vV6apmk7TdMwCAIMRgCXqaqqKvr9fpLneRqGYRYEQcnMhfd+Oh6Px9PpdGytHTnnRiLSUkq1RCQWkUhEQqXUlIgCrXUeBIGaTqel1rra2dnh58+fu+Fw6L/66qvV8Uw2wnA4lK+//tqHYejKsqyUUrn33kRRNGbmwBiTaq073vvxbDabnJycTIkods5xkiRhEAQKAQjcpnn6SavVXXUrkDr8WH+FucyDiPNX0r9FKVY0A431FXyXzHGD9a5Us/EV3RCdq9S/qByracAF09YZxtrJ1odDy+W7Yj288siaw+zZc9/YzxdcuXvVMPeL68ov2IfSeC4vWtLyOs7vg/Mh1co+aMzCRLSafCwFF0u1gaczLg9+vrIKaq57TbkuzvKucMnzclHrpisWfGHod+0yrSxv/cvxJ1uq7L1Bue7yCcOiZcelx5Lzx9bLybo/F5ehnuqCYOTc/Ivn9/LXVv2ZcZ3QY93pzfngphE0NJd50THkButanlEu3varS7lcrnULuCzgoEuyAFn+Z+ktesnnwrXfiuuuDWj8s9j7S7teFq/Ns+elGU7X3WY17qM6OKmPhTi1BQAAgM2HAOQDEBF+8eKFOjw81GmaBtbasKqqUERaRVG0RaTjnOt677ve+573vuec6zvn+kmSDKIo6j948KC/s7PTSdM0FRFDREEYhmG32w2TJNFKKZydwqWMMSpN0+Dhw4etdrtt8jxPtdZORMrJZDL7/vvv06qqktlsFltrk6qqEq11S2vdUkq1lFItrfXEWjupgxBmnimliqqqyi+//LLqdDqOiNy67rs2weHhoezv73uttdVal9bavCzLqdY6DIJgIiKj2Wx28uc///l4Mpm0B4OB2dnZoQcPHrDWOlRKXb0SgPdstcKC1ekYH6v9qjevSr+8BcRPLlFjvTeY64ZXqHOzVvg6FbxXXa197qr9a1RSXzrJNbbn0rym8eAF9ZoXV6XJ0s1mi5XL/NR6LxFP9VgvzSuxb6LZrdhSW5EbLmptnnFBK6F30xLk6vXflvdVlo370L+OutupS6e5Toy1MgOdvV+vnK9u5bA64bVa0Kx/tNn64VqjotzgPXE21tJbvtKusy65eCyPNRM3fq93o7JetKDVVEKus2dvEIA0VrIuACE6C+yWHqpbejLTouus+TkBN6ZZXRzCDwAAALhPEIC8f/zixQv1/fffmzRNTZIksfc+qaqqJSLtqqp63vu+UqqvlOq3Wq0+EfVFpGet7SZJ0u/3+929vb3egwcPOr1eL6H5gOZKKR0EgQrDUCEAgatorTmOY6O1TjqdTuicE6WUt9a60WiUWWujPM8j51zLWtvWWneMMV1jzCQIgjEzn3jvT6qqOiGik6qqQmNMkCTJtCgKlWUZTyYT+7vf/Y6++eYbLyKb1iWWDIdDHg6H/u///u/t//7v//Lu7m5WVZVh5iAMw1FVVe0sy47zPO+Mx+NWURRBGIZma2sriuM4uO0NACCiswoOorOKj/n9tXpMpcs+OG7vzTtf8w0/1d71h+BNt/99BEY3X8EF867cfa2KQ755yHChG7c4aIRm81/rWmVc3q3UNa4Nl3m3Pes29B2/AZguawHyNgtr/P8WL9b38el8UaXsJjsbUPuqEOQtNlj8O6lgfptdzWsqvN+Ja7T8eGerWvy61pSXur0vUe9gHy0Vfnl5csFksubvuTAE4QcAAADcIwhA3rP5mB+6KAqjtY6894n3PmXmjoj0vPcDa+0gDMNBHMdb/X5/YIzpa627VVWlURR1ut1up9frdeZdXsXoZgfehjpFq12lVVXliCjo9/tqNpsZrXXsnGsppTrGmF4QBNMwDGfOueOyLI8mk0mrKIqoqipNRGo2m6lOp8N5nrO1tvjmm2/k6dOn9vnz56vfrzaBEJFPkoQ+//xz0lpLnueGiALn3JSIxkVRjPI8P5nNZu0gCFp7e3st772V93HJMMBPdVE3IdfuPmRznKuk/MAbt1H78ppnEe9mm5b6Z/mJi3ofe1lufA32W1sz6PfZjrnhFeg/oQusmwdSH7P3985evfIe3sK1XsdXT/QxPAtXnaYuHsXXTAAAALiHEIC8PzwcDvnRo0f66OjIaK2jIAjioijaSqmu935rHn7sWGt3Wq3WdqfT2X7y5Mlur9frRlHUds6FzByHYRgPBoMoiiI8X/DOKaU4SRKzs7OThGGoiqKIiaitlCq11pUxpgyCoMiy7Hg0Gr3+9ttv2865JM9z7b3XWmtVVRWLCIsIG2OoLEt69OgRDYdDNxwOiTbnu6UMh0MaDof+yy+/pL29PTk5OSlEJPPeT4lowswj7/2JMaYThmEnCIIeM7sNa+0CAABzHyS/vnQdN+tA6V20APkgn8r34VMRYREAAAAAwMZDhfp7UocfW1tb5n/+538ipVSstU6NMR1r7Za1dltEdrTWD7TWu61Wa6fb7W7v7OzsDgaDTpqmLe+9JiKtlNJRFJn5IMu3vWlwzyilOAxD3e/3oyRJjPc+JiKvlHLMvPg7m82OtdbtyWQSVFVlqqoiY4yy1ipmZmNODyfGGPnTn/5EW1tb9Otf/1qGw6HfxBBERNyLFy+EiMo8zwtjTKaUmiqlJkqpsTFmxMw9EcmstWVZlo6IvNaa52OB4M0KAACn3uf52139tLmr5QIAAAAAgI8KApD3g4lITadT8+bNmziKolZVVW3nXKcoim3v/Q4R7Wqt96Ioepgkye7Ozs727u7uoN/vD3q9XpqmaUREJCKLHq8QfsD7wMwUBIEyxqh6HIt1rRmUUrFzLhoMBpqZA2OMLorCWGtNnuc6iiJFRFprzURUjwYujx49cvOWIJsSgBARyfz95v7lX/7FpmlaMnNurZ157ydKqbGIjK2148lkMvnxxx+zsixbaZqqVqtlwjBUWuur1gEAAAAAAAAAAADvEQKQd4+fPXumiMgwc9Tv91vW2o5zrue973vvd6y1u1VVPej1env9fn/vwYMHuzs7O/3BYNBtt9txEASGmU8vIUfoAe/ffHxkbr7ezr3wwjCM2u12Z29vT5Ik0UmSqFevXpmTk5Mgz/NARJRSynjvVZIkOk1TevXqFW1tbZXfffedEJH/gNv0znz33Xeyu7vr2+22jaKosNbmzDxzzk1Go9HEez8ejUbjra2taG9vjx88eBBrrYN5EAQAAAAAAAAAAAC3BAHIu8XPnj1TBwcHOkmSoKqqmJnbSqmuiNTdXu0R0Z7W+kEURbu9Xm/34cOHOzs7O51ut9uK49gYY9SVawL4wJRSQRzHqdY6CMNQM7PKskxlWaa11lpExHuviIiKomDvvdQ/g8HAz7vC2rgQZH9/X46OjnwQBLYoilJEciLKrLWz4+PjydHR0eT7778fP3jwIBGRoNvtBmmaajprBXNv1AEZxnsHAAAAAAC4GWMMvkgBANwCBCDvBg+HQyYi9fr1a52mqWHmSGvd8t53yrLs1wOeB0GwmyTJbhAEu7u7u9vb29tbg8Gg0+12W+12O1JKMaHXZLiDlFJaKcXGmICIyFork8lEnHPMzFxVlauqiq21Mh8PxBljPBH5v/qrv3JhGLr5AONCmzMeCBERhWHoq6qyRFQRUeGcy733s9lsNsuybMrMU611tr293bLWWhEJbrvM74KILP0AAAAAAADAzSilRGst3m/c9YAAAPfCvbtC+RbwcDjkb7/9Vne73eBv//ZvQ2ZOtNbtPM97RVEMqqrayfN8r6qqB8aYB4PB4MHnn3++9/Of/3zn0aNH/U6n04rjONRaa2ZWjH6v4A7iU1opZcIwjFutVm9vb2/v8ePHj588efIkTdNPlFIPsyzby/N8J8uyLWttp6qq1snJSURE5tGjR/rrr79WtEEh3+HhoYzHY/HeuzzPq7IsC6XUzDk3s9ZOq6qaFUWRV1VVeu+tnLrtYr8X93W7AAAAAAAA3rV1Y2sCAMCHhxYgP1Edfjx+/FgbY4LpdBoZY5Kqqtoi0rXW9kVke/6z22q1dre2tnZ+9rOfbQ8Gg26n00mTJEG3V7BRlFKm1WolxhgdRZEKw1BlWVbmee5FxDvnxDlXlWVZKaWqOI7L0WhU/frXvyYikuFwyMPhkGhDWoJEUeTTNLV5nldEVCilchHJiChj5pyISqVUpbW2SimPE10AAAAAAADAd0MAgNuHSvefhl++fMlffPGFSpIkiKIo9N4nIpI657rzQc8HxphBmqY7u7u7Ozs7O9s7OztbW1tb3Xm3V2EQBHre9RXARlBKqSAIgjiOW2madrvd7mAwGOxtb28/2NnZeZCm6a7WelBVVY+I0iAI4jRNQyIyT5480V9++aWadxt35w2HQ/nuu+8W44B47ytrbUlEuVIqZ+Zca10EQVAqpZxSCu2aAQAAAAAAAAAA7gC0APmJDg4O+M2bN3pvb8947yOtdauqqg4R9ay1W9ba7TRNdwaDwc729vbu3t7eYHt7u9vpdOIkSQJjjL7tbQC4qXk3bdoYQ2EYxkmS+MFgsKu1piRJ6OTkxI1Go8xamzHzrCzLLAzDPIoi/80338iTJ09kf39fRIQ34YqYly9fymAwcIPBwGqty7IsC+dcoZTKlVKF1rrQWlfGGMvMsgnb9FNgMHQAAAAAAAAAANgECEB+gnrg8yRJ9HQ6DaIoisuyTEWkKyJ97/0WEW2HYbgzGAx2f/7zn+9ub29vtdvt1jz8QAsc2Hhaa5MkScLM20mS6DRNlVKqzPN8Oh6PZ9baCRFNoiiKiqLwSinfarXcs2fPNqWlhBwcHEgURd5777TWlplLrXVRlmVhjMmNMUUQBOX8MaQCAAAAAAAAAAAAdwACkJ9gf3+fp9OpOjo6CsqyjIuiSL33XREZBEGwkyTJXhRFD3Z3d3cfPnw42NnZ6fV6vTSO41AphcHO4V6Yv5aDVqulmdk75ypjzAkzH1dVNdZaT5xzWZ7n5byrN/nzn//s//CHP9CrV6+EiDzd8bFAvvrqK3n+/Ll89tlnbjqdWudcRUQlMxfMnCulMu99lmVZdnJyMjPGhNZajqJIaa2VUmqjw876UMXMaPUBAAAAAAAAAAAbY6Mr5W6TiPDR0ZGazWZGKRV47+OqqtKqqrpEtBXH8c7Ozs7ez372s73Hjx/v7uzs9NM0bcVxHBhjDAIQuC+YmZVS2hgTBEEQGWMSImpba7vOuZ5zbstau1VVVbeqqlQpFed5HpZlqZ8+fboRY4EwM718+VLSNPVpmjpmtlrrKgiCQmtdMHNWVdV0NBpNv//++8n3338/e/36dZHnuXPObWxi0DxE4XAFAAAAAAAAAACbBi1A3oKIMBFxGIZ6NpuZoigia23CzKlzrqe1HsRxvLu3t/fg0aNHD7e2tgZpmraTJAk3/UpwgMuIiLLWBtba2Frbds71RWTmvc+rqiq01l5ErPfeeu/d06dP7f7+vicipjveCuTg4ECOjo6kKAoXhqGz1lbOuSoMw9x7P5vNZtMffvhhNB6P0wcPHoSPHz9WYRgqY4wKggBj/QAAAAAAAAAAAHxgqIx/C8+fP+ff/e53Ok1TE8dx6L2PiahVVVWnLMuetXaLiLaiKOr3er1up9Npt1qt2BhjmBn7HO4tZmattYnjuNXtdrv9fn/QarW2mXmnLMtBnue9LMtSa20sIuE333xjDg8P9Qa0ApHhcChbW1tea+2rqnJEZOcDoOda66lzbjIajSZ/+ctfxq9fv56ORqOiqirrvb/TwQ4AAAAAAAAAAMB9hcr4GxIR3t/f5/F4rEejUVgURWyMaYlI21rbs9b2y7Lc8t5vMXM3DMM0juM4DMNQa63R7RXcZ0opHYZh2O12O7u7u4NHjx7tdrvdPWPMrrV2J8/zvrW2XRRFIiLhbDYL9vf3NRGpecuqu0wODw/FGOPLsnTz1h9lFEWzIAgm3vtxURTjk5OTyXQ6nRVFcdr/FQbNAAAAAAAAAAAAuBUIQG7o+fPn/PTpU/Xq1SujtQ6NMbH3vuWcazvnOvMxD3plWbarqkq892YDKnYB3gmttUqSJNzZ2Wk/fvx48Nlnn+0MBoOdIAh2iqIYeO+7ZVm2vfet2WwWR1EUEJHe399Xz58/v/Pvk+FwKFEU+SRJHDNbZi6ZOTfGzIwxU6XUVGs9U0rlWuuKmR0z+9suNwAAAAAAAAAAwMcIY4Dc0P7+Pv/+97/XYRgGeZ7HVVW1nHOp1rrdarW6ItJrtVq9TqfTCcMwVkqh1Qd8NJRSHASBUUqxUoqMMVRVVemcK0VkWlXVCREde+/HSqnZfOD0qqoq9+WXX3o6HQfkTreY+O677+TRo0euqiqbZVmptc5FZOq9nyilpkqpmdY6V0pVCD8AAAAAAAAAAABuDwKQGzo8POSnT59qZg6VUrFSqiUibaVUNwzDXrvd7rXb7d7Ozk670+nEQRAgAIGPBjMrrTVprbVSipiZyrKsRKQiomlRFG9ms1mnKIoTY8w0z/Oo3++XZVlWnU6HRYTu+NtFXr58KZ999pmfzWYuiqKKmQsimjnnpkVRTJm5DkBKrbVj5jsd6AAAAAAAAAAAANxXCEBuaH9/Xx0dHRnvfe035c8AACAASURBVGKtbTvnuszcC8OwNxgM+p988snWzs5Ov9/vdzudTitJEqO1vtM1ugDvAzPrKIqira2tXhzH1Ol0yuPj46PXr1+/LsvyuCiKaZIk06qqiu3t7eqHH36w826w7nRgcHBwIOPxWLrdrhuPx1UcxzkzT/M8n2itJ8w8nXeLVd6HLrBEZPEDAAAAAAAAAACwSRCAXJOI8IsXL9TR0ZEZjUZRq9VKrLXtsiy71tpeEAS9MAy7/X6/vbu7m3a73SRJksAYgxYg8FFSSrExxiRJkmitvda6a63tjMfjlJlbzJxYa2NjTH58fFxMJhO1v7+/Ee+VN2/eSFEUPkkSmyRJUZZlFobhrCiKWaMFCLrAAgAAAAAA+Mh578laS0phGF4AgNuAo+/VeDgcqhcvXigi0rPZLHTOxUVRpEVRdKqq6pVl2bPW9pi5G4Zhu9PpxJ1OJ4zjODDGKAQg8DGad4elwzCMklNpEAQpM7dEpOWcS7z3sfc+JCLT6/XU4eHhnX+vDIdDISK/s7PjgiCw3vsyDMOciDIRyYgoV0oVzFwHIPeq6QQOZwAAAAAAAAAAsCnQAuRyPBwO+dGjR3o6nWrvfUBECTOn0+m0673vF0UxqKpqEARBfx6IxNZaIyKoJQRoEBHlvQ+stbH3Ppn/xEQUaa2DOI7Vl19+edvFvJb9/X0hIj+bzdzu7m6VZVmhtc6JKBeRnJlLZrbM7O/DGCAIPQAAAAAAAG6GmcV7T/fhOyEAwCZDC5DLMRGp6XRqxuNxyMyx1rrlvW8757rW2i1mHkRRNIjjeBCGYZeZEzoNllBjCDAnIuy91865wDkXO+daIpKISGytjcqyDF69eqU7nc4mvG/k8PBQdnd3/e7urrPW2iAICmNMTqetP3LnXOGcK7IsK7Msq4qisNZa773f2BNfhCAAAAAAAADXJyIIPwAA7gAEIBfjZ8+e8evXr3VVVUYpFWRZFltrW0SUlmXZdc71giDo93q9/vb2dq/X63WTJIm11poQgAAsMDOJCDvnAmttbK2NnXOx9z4SkdBaGyRJov7jP/5D0Qa8d4bDIf3zP/+zfP/9977X61ljTFUUReWcK4morKqqmEwmxfHxcXF8fFyOx+Oqqiq3yQEI0fKA6BgYHQAAAAAAAAAA7jp0gXWJra0t9fnnn6uiKExVVaH3PrHWpmVZdqqq6sRx3G23290nT5709/b2+nt7e+3BYBCdjvmsb7v4AHeGiLCIKOecmbcCibz3ERGFSqlARLQxhn/5y1/WV8ncdpGvIgcHB/Q3f/M37g9/+AOnaWpns1lFRKVzrjw+Pi6YOZtMJuPt7e30wYMH0cOHD+NOp8PGGATPAAAAAAAAAAAAHwACkAsMh0MmIh6NRjoMQ5PneaS1bllr06IoOtbaDjN3oijq7OzsdB4/ftze3t5OkyQxYRhi4HOAFd575b033vtQREIRiZxzofc+iKJIl2WpkiTZlPeNfPXVV0RE/ne/+507PDy0SilbVZVl5moymRR5nmc//vjjdDKZTEUk7XQ6ptVq4ZgLAAAAAAA/Wd0aG62yAQAALofKuAu8fPmSDw4OFBEZ732olIqJKLXWdp1zvbIsu9bajlKqnaZp2uv1kn6/H2mtkX0ArKhbgNTjgFhrI2YORSSqqioIgsBYa9VkMuHnz5/Xb6A7fSbPzCIi9M0333jnnMuyzFprK+99lWVZ6b3PnXMzZs663W6R53ninLvT2wQAAAAAAJsD4QcAAMDV0BXLBQ4ODpiIVFEUOs/zUETioig6ZVl2y7LslWXZKcsyLcsyds4ZpZTSWtM8/ah/AOAMi4j23gciEjjnQudcwMymLEttrd3I49GzZ88kTVNfFIVzzjnvvXPO2flP5ZyzImKZ2dMdD3UusyFdkwEAAAAA3HsIPgAAAK5vIyscPyAVRZF2zgVVVcXe+5SIOszcNcZ0tNYpMyfMHHjvtYigdhDgAiLC3nvtvTcisvipqsoQkTbG8AZ1gUVEp61AiEh2d3c9EXkR8d575713ImKJyCqlrFLKbXIAgi9YAAAAAAAAAACwiRCAXGI2m/F0OlVEZKqqCq21CTOn7Xa7vbOz09nb22vv7Oy04jiOMLAxwMXmXWDxfBwQ7ZwL6iCEiLT3XhVFwUdHRzwfW2NjMLO8evVKRMQTkXfOOWZ2zOyIyImIIyJ/y8UEAAAAAIB7hJnRQhsAAOAaMAbIBb799luOooiTJFHee83MgbU2StO01el02oPBoLe9vd0bDAbd7e3tOI5jg5MPgEuxiCgR0SKi6XR8HeOc09Za7b1XDx48oBcvXrCIyCa9n168eEG/+MUvqA5BmNk559y86yunlPLz1iIAAAAAAAAAAADwgSAAuURRFGyM4TAMlXPOiEgQhmHY7XaTTz75JN3b22v3er00SRKjlFLWWtJaS+NKjM2pwQV4jxrvByUimpn1vNs4TUSamVlrzScnJxv5njk4OJDj42Px3ouIeBHx8xYgvvEjCEEAAAAAAAA+Lt57EhESEYrj+LaLAwDw0UEAcoGjoyP+5JNPmJlVURRaKaWVUsY5FzjnAmutKYpCT6dTNZvNWGtNURRRmqbUarUoDEM0RwVY4b1ftACZD4iu6TQUUdZazvOcO53ObRfzrcxmM0nTVLz34r33ROSVUnUIIrSh4380YSwQAAAAAAAAAADYJAhArmCt5SAIWESU997MZjN9dHTExhg/Go2qIAgq770opUyn0+HHjx/z3t4ea63JGOxegFo9Dkg9Fsg8BFHz95ZSSvHOzg4VRXHbRX1r1lohIlFK+bolCM1bgDCz3IcA4T5sAwAAAAAAAAAAfBxQQ3+F0/GMWdHpgPF6MpmoyWRCf/nLX0pmzokos9bGURTxgwcPlLWWkyShNE1vueQAd8dq+EGn7yellFIiopRSzPMmU8+ePbvdwv5EzFx3hSXOOaF7FH4AAAAAAADA9eF7IADA7UMAcg3eexYRxcyqLEsuy1KKonBFUVRVVZXee5MkSeCco08++YSKoqDTHnAAoOl0bHNmmgcg85YgyjnHxhgaj8f8r//6r/yb3/zmtot6Y1EUibVWtNbivRead4HFzIsWIBgDBAAAAAAAAAAA4MNBAHKJoihYRFgpVV/Brqy1XJYlj8djmU6nvqoq772XsixlMplQnufknEPKD7AGM7P3Xnnv1TwI4ZrWejFozvPnz5k2cMwMrbWcNmoRIaLFX6LTliG3WzoAAAAAAAAAAICPCwKQa3LOETPTvAsf8t4zETHRaZPG+gcA1pv3cLUIPRqtQe4dEalbgRDdkwHQAQAAAAAAAAAANo267QJsgnnYUd8mmgcfzccQfgBcTkTq981S+DEPFe9NEDIf94O896dNQDb82FBnVKvbUf+/6dsHAAAAAADwrqELZACAuwMByCXKsmRr7YUVs/OKv42v4AT4UOoQpK5UZ2ZW6vQwVFUVT6fTexGEeO/vzclufXxb11gHxz4AAAAAAIBlze+C9+V7IQDAJkMA8naaXdsQM6+tHAQAuE8QeAAAAAAAAAAAwCZBAHKJMAzFGLOU3DeaMQpCD4Cbqd87dUX6fDwdIiIKgkDSNL0XNexKKW50+XVv4RgIAAAAAAAAAAB3GQKQS0RRJFprUUrJmvBDmFmUUs2A5BZLC3C3rTYDltOBQM69jzZdHXwopU5He79Hx4X7tC0AAAAAAAAAAHD/IQC5BqWUzH+8UsrN//q6Qrc5uBUqCAEuthIk3lve+2YLEJ7/bKTGeC23XBIAAAAAAAAAAICbMbddgLtOay3OOWmEHosfrbVEUSRhGEq326WtrS1qtVpkjEFlIcAFmq2oalrrexGIOOc4CAIqy5JEhOuf2y4XAAAAAAAAAADAxwgByCWOj48pDEOK47jupqcOQZxSyodh6JVSvtfr0c7ODj169Ij6/T7FcUxKoXENwEXmrUB83bqKiMg5t9EhSFEUrLUm7z0rpZiZyTlXd4GFIAQAAAAAAOAj5Jwj7z1prW+7KAAAHyUEIBfY2toSIhJjzFL3V1prq5RyzOzjOJZOp0O/+MUv6NNPP+UnT57w48ePqd1u44MNYI06SJyPgi5E5JVS9Xggt128n8wYw845Vkqx977u+mrzNwwAAAAAAAAAAGADoZnCFeZd89StPiwzW611pbW2SZK4ra0t/+mnn9Kvf/1r/tWvfsV7e3vcarXQAgSgoTHuhyciqbuTq7vAUkpJEASLFiBfffXVxrYG0Vqz956994pOj7GK5i1A0AoEAAAAAADexn24YOxjVfd6AAAAtwMtQK5QVZVEUeSVUpaIKq11qZSqlFI2DEOXpqns7u7Kw4cPaW9vj7XWOCsBWENEFl1f0WmoKFrrRRBCRNTpdOQ3v/nNxp4czscAqcMORURKRNT8NuNLCwAAAAAA/BT4TrGZ7su4lwAAmwjNFC4RRZHEcey11k5rbYMgKI0xpda6MMaUxhhrjLHzq9nxYQZwiXrwcyLyWmunlLIi4uou5bTWvtvtyosXL267qDf28uVLbrVabIxh7z0zsyIiVf+tA5BbLiYAAAAAAGw4EVn8wN3V6AUBAABuGVqAXODx48dCRL4sSy8izhhjtdaFtTY3xhRa69IYUxljnNbaK6XuxRgGAO+RKKW81toxsyMiZ4yx88HQvfdeyrLc2BPEoihYKcVaa2WtrYMPTfMusJiZ0AUWAAAAAADAx6MOQkSEmt0+AwDAh4MWIJdI01Ta7baPosgGQVBqrXOlVG6MyYwxxbxFiJ1344N0H+AS8y6vXD2ejlLKaq0tEbkgCFwYhhv7/nn27BmVZcnMrJxzioh080dENMIPAAAAAACAjxPGAQEAuD0IQC7w8uVLmU6nUpali6LIaq0rY0weRVEWBMHMGJMbY8ogCKp5pS4+zAAutuj+ak34YZ1zvqoqX5alHB4eblprKj48POQ4jtkYw8YYxcxaRHT9l05bg2zURgEAAAAAAMDbQz0RAMDdgC6wLudpXmEbBEFJRLm1dmaMmQVBkAVBkM9bgSAAAbhCPQC6Uqoe/8MysyUip5Ty1lr58ccfb7uYN8VERN9++y13Oh323isRUUopbYwxRBREURQYYzQzK4yCDgAAAAAA7xK+YtxtaPkBAHD70ALkAgcHB/L69WtJksRFUVR57wul1EwpNQ2CYGKMmYRhmIVhWGitrVLK33aZAe6yugssY4xVSlVKqYqZq7olSBzHsrW1tUknh0xENBwO+YsvvlDWWq211sxs2u120O/3o0ePHsW7u7txr9eLwjA0SikccwEAAAAA4NqYeRFyNMOO5v2rjwEAAMAZVMZdYDgcSlEUPssy572vjDF5EASTIAhGxpiTOI5HcRyPoyiazUMQd9tlBrir6jFytNZWa10aYwqlVBEEQcnMlTHGGmM2LkQcDof85ZdfqiiK9NbWlmZmQ0RBv9+PPv3009Zf//Vf9371q191P/nkk7TT6QRBEGz8MRdfrAAAAAAAbo+IEDOTiCx+AAAA4GIbXxn3Pv33f/+3DAYDV1VV5b0vwjCcaa3rEGQURdEkDMOpUqoQkcp770TEy+kZCM5CABqY2dcBCDOXWutCa13OW4K4siz97u7uxrxvRIT29/d5b29PGWO0iBgRCUQk6HQ60cOHD1tPnz7tfPrpp529vb1WmqaBMQbHXAAAAAAAuLFm2IHQ4+5DOAUAcHegMu5i8pvf/MZHUeSzLHPW2sp7nxtjZkQ0jaJorJQaEdFJWZYnWZaNZrPZtCzLYh6E3Hb5Ae6Mxvgf1hhTGmNyY0xBRKXWugrD0G5vb/ssy+Srr77ahACRX7x4oQ4PD/W///u/GxEJ0jQNgiAImTkMwzBqtVpxv99Per1e3Ol0wjAMtVLq3jSfWG1yDwAAAAAA715dt4Bz783RrA/yfuM6OgAAuHcQgFziq6++kq2tLT8YDJzW2sZxXFprc6XUzBgzYeaTqqqO3rx58/qHH354/ebNmzfT6XRqra0ECQjAEqWUn4+XUxpjCmYutNZFGIZlFEW2KAr/2WefbcT7Zjgc8u7uLne7XZ2mqSmKIlRKRVrrSCkVMXMUBEEQhmEQhqE2xmil1L0YBL1ucr96GwAAAAAA3o/VEKTZBRZsBDxRAAC3yNx2Ae6y+cmF/Pa3v/VffPGF1VpTq9UqyrLMnHMT59zJaDR6Y61tHR8fB5PJRD958oSDIAiMMQEhYAIgonMtQIogCHIRybXWhVKqJCJrrZUsy4SZ7/zJ4f7+Pv/bv/2b2t3d1cfHx0EQBKH3Piai2BgTi0jonAu894rmg6UDAAAAAAD8VHX4gQuRAAAArgcByOWEiOjx48fuzZs3QkTknCvb7XaWZdlERI6rqoqOjo7CLMuMiIRhGAZEFHU6HZMkicyv/ub7cOU3wE2IiHfOibXWlWVZzGazLM/zmYjMRGSmtc601vl8TBBrjHHj8fjOhx9ExIeHh9ztdnVZlsYYE5Vl2fLet5i5JSIt733svQ+ISInIRr33rbVUVRVVVUWj0Yim0ylZa8k5d9tFAwAAAAD46KHlBwAAwM0gALmaDIdDIiI/HA7p6dOnlbW2MMbMRGRUlmWY53lUlmWklEqDIEittWmv1wu2trao3++HSimttd6oSlCAn8p7L9ZaN51Oi+l0OptOp5PJZDKtqmrKzBkRZVrr3FpbGmNsp9Pxf/d3f3fnz+SHwyETkXLOKWY2cRyHVVUlItISkdR733LOxd77UEQ2qgWIiFBVVZRlGY1GIzo5OaHRaER5niMAAQAAAAC4I5pdYWFsvrvJe4/xPwAA7ggEINcjRETD4dD/4z/+ox0MBkUYhtMsyyLvvdFaRyISj0ajTlmWnaOjo3R7ezssy1JFUaTDMFRa69veBoAPynsvRVHY4+Pj7M2bN+OTk5OToijG1tqptXYWBEEmIrkxpux0OlWn0/G0IX2jDgYDJiLtnAustbFzruWcS0UkZeaW9z6x1obee71JLUDqAGQ0GtFf/vIXOj4+ptlsRmVZkvceX6wAAAAAAO4InJtvBoQgAAC3DwHI9QkRyZs3b1wURbbT6eRBEEydc2FZlq2iKFplWR7PZrNelmVdZk62trZCa20sItjP8FHw3kvd8iPLsnIymeQnJyfj4+Pjk5OTkxMRGRHRVCk101rnSqnSe1/NZjOntd6EAIT39/f5T3/6k4rjWHvvg7Iso7IsU+dce94CJPXexyKykQGIc47yPKfxeEzj8ZjyPF80s6+b2te3mRnBCAAAAADALcF5+N01Hwfzrn+/BQD4KKBi/ub81taWjaKoYOasKIpARGLvfVIUxXFVVb2qqjrtdrtVVVVCRG0iCm+70AAfgvdeyrK0k8mkGo1Gs/F4PDk+Pj4ej8dHWZYdKaVOgiAYh2E4DcMwY+bCOVcZY+wPP/zg9/f3b3sTrnR0dKRGo5HO89wwc6iUSqy17aqqut77jve+7ZxLnHOh917ThnWB5b0nay3leU55nlNZlqSUWny5avY3jL6HAQAAAAAALoYQBADg9qnbLsCmGQ6HQkSuKApblmWhtc689zNmnhhjxlrrkTFmHIbhJAiCnJkdPvDgY+Gc81mW2R9//DH79ttvx3/84x9PTk5Ojr33R1EUHRljRlrriTFmFoZhbowp2+121ev13KtXr2QDrmDi//qv/1JZlumyLIPZbBZlWdaat/poO+faRNRyziXW2lBENqoFyDrNVh8AAAAAAABwM6gTAgC4XWgBcnNyeHgo+/v77uTkpNJaFyKSicjUez9WSp0YY46YOXXOtfM8785mM50kiWitjVJK8QbU8gK8DRHx1lo7nU6z4+PjydHR0XEYhkda/3/27mQ3kiu7H/85d4g5h8gkWUVJthqCWzZYbgOGjAYM2FAZaBjwA/AV7J1fQVmvob034taAt+q1oZUgon+N/gvqbrmqJBaZzCmmO5z/gplUFkVWcU6SdT4AkWQyM6aMiLxxv3HvlQdSykMhxFhKORNCHLf+GI1GTinld3d3Ce54F1jb29uolBJxHEtjjBZCBNbaCAAyrXUWBEELEVvtdjtJ0zSUUkpEvFdB83JXVwBHzeqJCIQQHIYwxhhjjDG2IifL4FwmZ4wxxs7nXlXM3RWLViDWWlPXdeO9L+eVuhOt9aFSaui9P6iq6mAymQwnk8l4Op2W1lpDRDwCFnuwvPfknLN1XVdFUUym0+morushIg6jKBpqrcdSyhkRVVLKOssy8/z5c/ff//3fND+u7jJ88uQJvvfeewIAlNZae+9DIoqJKFVKtTqdTmtzc7O9sbGRtdvtOAxDJYS414HnaaEHZ7iMMcYYY4ytzmI8Pg5B7rbF57PoZpgxxthqcAByObS9ve3TNLXj8biRUlZENAuCYCSlPCCiH4uiePn8+fPnf/jDH/7v22+//WFvb29YlmXtnOMAhD1YQggvhLBa6zIIgolSaqi13tdav9Ja7wdBMIqiaJplWRmGYaOUsr/61a8cANz54+KLL74QvV5POudUHMcKAAJEjIwxiXMui+O4/fjx4+7f/M3f9H75y192PvjggzTLskBrfa/Os8vhxqLAftrFFYcgjDHGGGOMrQaXxe8HRCTv7/ylLmOMPXjcBdYlISJ98cUX/sWLF1Yp1UgpS0Sc1nUdCiG0MUYdHh6qqqq0MUYopWQcxyEiyjiOQQghhRB43+8OZ4yOeOecr+u6sdaWADBDxMk8FDwUQgy11odCiAkillrrmojMjz/+6KbTqZ+3/rizty8REX755ZcIAGI8HsvDw0MthNDe+9A5FwNAEgRB0mq10vX19XRtbS1OkiQMgkAIIe5VAHKaxR1mfJcZY4wxxhhjq7EIPd5UHuey+t0jhCAAACkl1XUNxhh47733aG9vb9WLxhhj7wwOQK5gd3eXnj9/7uI4NkKIWik1i6JIe+9l0zSyrms1Ho9D730QhmGYJEkCAMo5h0mSaKXUve8ehzHvvbfWurIsTVEU5XQ6nRljpog4VkqNEPEwCIJhHMeHWuvJZDIpkyRpmqaxf/7zn/1//Md/3OnwYw5brRbu7e1JY4wyxmgACIgoJKLIex8DQBKGYdxut6Msy8IoivSqF/qyFhdXy3eW8V1mjDHGGGOMrd7ipqTFTUoLHH7cXYhIRARaawrDkL777jtI03TVi8UYY+8MDkCuYDAY0BdffOG///57i4gNAJSLlh1EJBBRW2sTY0x0cHAQee+joihEv9+H9fX1NMsyBO6GjN1zzjlflqXZ39+fjsfjw8lkMpzNZofe+0Ol1EhrfUhEIwAYl2VZtFqtSkppfvzxR5fnuYc7Hn4QEe7s7ODf//3fiyzLxGQyUVEUaWNMQEShtTZSSkXW2tAYo7339/qYXr5wOusiii+uGGOMMcYYWx0uj999QghCRAI4GgOEbyhjjLHV4QDkamh3d5cAwKVpatI0RSklSCnJWouTySQgoqRpmvDg4CCYTqe6aRq01kIYhoumkCiOcHdY7N5Y6vaKyrJsptNpcXBwcDgcDofj8XgfAPaJaCilPJRSHiqlRlLKqda6zLKsllKaOI7dv/3bv935AAQAYH19HX/3u9/JsiyVtVZ57wMiihAxIqLIWhtZa0PnnPbeCyK618fyaRdUZ40HwgV5xhhjjDHGVmPREoQDkbtp3krnuAss/pwYY2w1OAC5Hj4MQ5tlGUgpF+m+1FpHQoikqqqwrutgPB5rRFRBEIgsyyQAIBGJKIq01lpyAMLuC++9N8a4uq7tdDotR6PR9PDwcDQajQ4mk8m+1noYhuFhEAQjpdQEAGZCiDLLsvqv//qvmy+//NI9ffrULwqDd12r1UIAEMPhUAGAJqJACBESUQgA4XwskMA5px5CALJwMtw42TUWF+AZY4wxxhhbDb4R6W5bDH4+rx8iYwwoxVVwjDG2Cnz2vaLBYEDb29v0m9/8xjvnXBRFBgCwKIpSCDEhokhrrQBAEBE2TYPD4dAjIhVFYaqq8vPusEKl1L3uOoe9O6y1fjabNcPhsByPx+PRaHRYluW+c+6VUuqVUmpfKTXUWo+UUrMwDCsAMNPp1O3u7tLTp0/vw7gfAADw7Nkz3NraQgCQxhglhAgAIASAiIhi731IRAERKe+9vM/hx2Kg87OCDw48GGOMMcYYW53lVtkLHITcPcs3+i0GQWeMMbY6HIBcHX3xxRd+Z2cHhsMhAAB479F7X4VhOLXWBs45qZQSRITWWhyNRlQUBZRl6YkI4zhGpRRKKVEIIXBuxevF2GvoJ76qKjOdTsuDg4PxcDg8nEwm+9baV0T0Sim1r7U+kFIeIuJECFEYYxqttU2SxH3//fd+a2uL7kvrDwCALMvw+fPnEgB00zShlDJCxFgpFUdRFANAFARBoLVWiCge0uG76PLqZDDCYQhjjDHGGGO347RuaE+Wzx/SNchDgIjH17zc9xVjjK0WByDXABGJiI5DkCAIoNVq4Ww2k4iolFKLAbC8MYbqunbOOee9t0EQUJqmhIiOiLIoigKttZJSylWvF2PLvPfOWmurqrKz2Ww2Go3Gw+HwcDQa7c9ms1dSyh+01ntBEOwJIfaVUodBEIyFEIUQov6///s/G8ex++1vf+vnLUDuha2tLfzd734n4jhWiBg456KmaRJETNM0TbMsy7TW6cbGRtxut4MwDMVD7c5uEYQwxhhjjDHGbsdpIcfJ+vSTXdUyxhhj7CccgFyTebLvB4MBbW5uQtM0NsuyqigKKaXEuq5x/jqs65oAgKy1bjwe+xcvXtimaZqqquza2lo7TdOYAxB211hr3Ww2q4bD4Ww8Ho8PDw+HVVUNnXP7UspXUsq9+eNrrT+EEHXTNGYRfgwGAxoMBvcmANnd3cX19XUJAHreoisiokRrnaZp2srzvJXneavb7WZra2tRkiRKSnmvrzzedEHFNy8xxhhjjDF2d3DocXfNB6jnCyjGGFsxDkCuFw0GAxgMBm5zcxOcc9jpjcEVbQAAIABJREFUdHA0GkGaplQUhQcACMPQSym9c86Ox2PfNI2pqsoYY3wURVJrLZRSEpesesXYO2lRViMiorqum+l0WhwcHAyHw+FwMpnsG2MOAGBfKbUvpdyLomhfSjmMomgkpZxIKQshRP3111/bg4MDPw8+7lMBEAFATCYTmWWZAoDQORc75xJEzOI4bm1sbLTef//9VrvdTrIsC6Mokg+xBcjJEITL8YwxxhhjjK3WWWP4sbth0QXWfBwQ0lrzRRRjjK0AByDXjwaDARER7OzsmKqqoNPpQFmWlGWZr+sayrL0QohFd0K+KAqLiF5rTb1eTwVBAIgIQRBopZRCRP6c2EoQkbPWOmutqapqMpvNDieTyf5kMtmfzWZ78/E+9qWUB4j4ChEPwzAcOeemzrnCOVfHcWweP35s//M//9Oven0uAQFABEEgnXOBtTYyxiTW2lRKmWmt0yRJkjzPo3a7HQZBoBERhRCrXu4r44soxhhjjDHG7q7TxgDhMjxjjDH2c1yxfkMQ0ROR/eqrr+jFixektfaHh4cOEX0cx8Y5V9V1XTnnaiKqjTFmMpm4H3/8EeeVzbbb7WZJkqRBEPDnxG4dEZG11pZlWU6n09lkMjkYj8f7VVXtAcCe1vrHIAj2lFIHQRAMhRCHUsoJAMziOC6FEJUxxgCA3d7evm/hBwIAPn36VKRpKoUQumma0HsfN02TWWtbSqmWtTYDgFgIoeWR+598wE/hhxCCL6IYY4wxxhi7w7gVyN1EROC9P24FwhhjbHW4Yv0GzUMQ+PzzzyHPc+r1em5/f98BQENEVRiGTVVVzjnnEZGqqqKXL19CVVWuaRqvlAJ1RBLRoicsPJr0cQGHSznsqmipS6PjLqq8994YUxdFMR0Ohwej0WivKIpX3vtXSqk9pdQPYRj+qJQaJklyCAAT51yBiFW73W6UUuabb75x29vb/p4V+o7Dj1/96ldyNpvpOI61MSYiopiIUillJoRoAUBKRBERKXhAx+Li/LLo5urkoIrc/RVjjDHGGGOrx+HH3YaIi2ttUkqRc47a7TYdHh6uetEYY+ydwgHIDUNEPxgM4OOPP6avv/7aP378mADASSktEfnxeIzGGAQAMMb4yWTihRBGKWWyLPNKKee9b5xzkoiUlFIGQaC01lJKKbigw66KiMA5540xzjlnnXMOER0imqqqpkVRDCeTyd50Ov2xrut9ANiXUr5SSu0lSbIfhuEhIk6SJCmstXVZlrUxxv7d3/2de/Lkyb0b82MwGODz58/le++9J+M41tba0DmXAEBCRFkcx60gCLpZlnXyPG/HcRxLKdVDHKvnAa4SY4wxxhhj9xqPyXf3ISItbgJcPFprQSmugmOMsVXgs+8tGAwGnohob2+PsiwDKSUFQeDH4zFGUSSJSBhjyHtvjTFmNpvVSqn64OCgcc5VWuuOtTYEgDAIgrjb7UZpmkZRFPEA6ezKFl1dTafTejabVcaYGhFrKWXpnBtPp9P9qqr2jDF7zrkDpdRQKXUQhuF+GIaHcRxP0jSdIWIdBEHzww8/2E8++cTBUmuSewSfP38u0zRVAKCdc6EQIvXeZ03TtMIwbCdJ0un3+3m/3+91u91up9NJgyB4kAHIafhCizHGGGOMsdu33NJjucU2twK5e5aumch7D0REUkoCABgOh/Do0SOaTqerW0DGGHvHcABySxCRBoMBffrpp64sS5hOp7S3tyeiKBJCCFBKOQCovfeVtbaYzWazly9fFq9evZoiYl7XdSqEaHW73TYRdZRSKgxDuer1Yvef956qqrKj0ajY29ubzGazCRFNgyAYI+LIWntQ1/UrInqltT5ExBEijqWUh0Q0EUKUiFjHcWyGw6FbhB/3rNsrAADc3t7GMAzF48ePlXMuDIIgIaLMWtsmog4RdbMsy99///3eo0eP1trtdp6maRxFkZJS8hUHY4wxxhhj7MacvBmJQ487jZZbgpy0vb19366XGWPs3uIA5BYNBgMaDAYeAGBra4uCIKgPDw9RSklRFDnvfSOlbOYDpJd1XVdEVHrvJ3Vdt7XWHWNMnaapDYLAeu9jIYQCAIGIUmstgyCQUkohhOCSEHuNn5t3deWstR4RyXtvZrNZcXh4ODo4OBhNp9NDABiHYThUSh0i4gEi7iulhs65iVJqAgAza+1UKVXWdV13u91mOBy6ra2t+xp+AADAkydPEABkWZY6juOwaZpUCNFumqZjre0EQdAWQrTjOG612+200+nEWutQSvkgW2MtmtYv7ixbPMcYY4wxxhi7HctlcYCj0GPequC1n+X/s1tH1lqy1npjjJtOp81kMjFVVTljjJ/3ugDee4iiCP7whz/As2fPVr3MjDH2zuAA5HbRYDCAeQhCURQBAMB0OvVN0/ggCAwAGCJqmqZp5pXU1jlXNU1TaK0rpZTZ3983QohmOp2miBgQkQrDMMiyLGy322EYhpoDEHaS957qunbT6bQqiqJumsbMx6JpiqKYTSaTw6IoDsuyPASAQ+/9UGs9DIJgKKUcCiFGYRhOhRCFc64UQpSj0ajpdrvmhx9+sN9++63f2dmhwWBwL2vIB4MBAoAoikJ2Oh3dNE2IiIkxpmWt7Tjn2vOfTAgRa63DIAi0UurBtcQiouOLqpOWm9p774+fY4wxxhhjjN2808IOLo+vFhGBtdZPp1MzGo2a6XRazmazejKZHAcgSimSUtJwOFz14jLG2DuHA5DbR4PBgIgId3Z2IIoiKMuSAMCHYWi01tY5Z5xzVinlhRDOOdcAQAUAVVVV9d7eXjWdTgspZeq9jxEx6nQ6yaNHjzKttdRaSwAQq11Ndtc453xZlmZ/f3/26tWr6Xg8LpVStRCics5N67oeOedGQoiRlPJQaz3UWh8qpUZBEBxKKSdSyqKu61pKWQNA/ctf/tJ8//337h//8R/9J598cm9bfgAAfPPNN/jkyRORJIk0xmghRERE6Tz06Djn2tbazFqbWGtDInqwx9jiourk3WTe+5/dfcYYY4wxxhi7Ocshx+JGpOXyOls9OrqL1Y1Go/pPf/pTMRqNZlVVlURkiMgLIcgYA845SNOU6rpe9SIzxtg7hQOQFZlXFPvBYECbm5sUBIGfjwPinXPeGOMBwBORA4BaSlkSUWGMKcfj8Ww2m00QMfPeJ0KI1FrbiuO47na7TikVG2O0917Mu8OSSik576bnwVbasiNE5J1z3jnnvfeeiDwi+qZp6qqqyul0enh4eDgajUZTKWUphCiEEBMiGnvvJ0qpsdZ6pJQ6DIJgHATBREo5UUoVQojKe9/s7e3ZLMvMX/3VX9n/+q//on/5l3/xq17vq5p3fyUAQM0Djth731JKdYIgyKMo6rXb7bzb7bajKIqklAoAHlwCcDL8WA5BTl58nfXedxGHQavxLu9zjLF3E3/fMPZmD61scFo3tItW2EopiOMYAAA6nQ5kWQZBEIAQfMl/2xYtQMqytKPRqN7f36+bpmnCMLRKKa8UV70xxtgq8Vl4tRatQWhnZ8d/9NFH7ttvv3VSSieEMN57E4ZhjYhTABgTUatpmlFd123vfct73wKADBHbSqnOaDSajUaj0hiTKaVC773SWgdhGEZZloX6yKrXmd0w55yvqsoWRdEYYxrnnFFKNcaYsizLaVEUh3VdD6uqGgshpkKIaRAEYyHENIqiCQBMpZQTrfVESjkDgEJKWc5mszoMwwYA7Hxf9YjoAeDeX2UQET579uy4+6u6rkPvfeKca2ut8yRJ1nq93nqe52sbGxvdLMtSKaV+aON+LIcf3vvjH0Q8vpA62QJk+S60y26Oh3ahym7PWWEce/ge2On3wni/Z4yxd8PJsfiWz/9KKWi325DnOeR5Duvr65AkCUj54HrovRecczQf/8NMp1NT17UVQjghhBdCEACQlJL4O5wxxm4fByB3wHJrkE8//ZS+/vprH4ahyfO8qaqqBIBQaz0holEcx5kxJpuHH23nXBsRO0qpcVEU4x9++GGslMoAIHHORUmSpN1utyWEwFarJQCAS0MPnHPOF0XRvHr1ajabzYqqqoowDGeIOPPeT5xzh2EYHnY6nZGUcqyUGiulRlLK2TzwmAkhCmNMEQRBVdd1I6VsxuOxAwC3u7vrYb6/wgMIPwAAnz17hgAgkiSR4/FYe+8j733qvW8LIXppmq598MEH648fP17v9/u9LMuiKIoe7Fg73ntwzh0HIUKI48ezmuBfpSL6Te+9SrDCHj6+gLwZt7Fdr3Jc8znh8uHfbR8z/FldP/5eZOzhO9nq47RHRIQwDF8LQDqdDrRaLQiCYDULzo7NPyOapx1ERCSlJOcctFotCoKADg4OVr2YjDH2zuAA5O6gwWAAROR++9vfegBweZ7bPM9NWZa1tbYhoso5VyVJUgDAzBgzM8bMiKgQQkybppkcHByMASAjosQ5l7Tb7UxK2Wm1WpVSKhFCBES0uGo6+bjsteeW3vPTC5Yuvk77/2Vfe1MuO9/bGtdiqZuhN87vxP9/9ntd13VRFOV4PJ6Mx+NpWZbTIAgmSqkpIk6IaBxF0WEcx2MhxCgIgokQYqyUKrTWhbW2klJWZVlW1loThqFttVpub2/P7+7u0meffXavx/o4aTAY4Keffir+/Oc/y++//17XdR157+P5MZQBQFtK2cmyrN3tdtt5nqdaa6WUEvDAusBatPTQWkOSJFDX9Wt3mi0CkcVrF8+dvBvtMt70/rP+d1YF0HmX5TorkBbb5bzexcqrm6p4ve1tedH1OO/ycZjD2+Ci3rS97so5ZhWf6UXX/arLuIpz0FWW+a7sG2x13rVz7X3c509+Rqd1USuEACklJEkCa2tr0Ov1IE1TCIKAW4Cs2PxamYiIEJEQkYQQZK2FIAjerQOQMcbuCA5A7haaF9AIADwAwGAwsJubmyaOY9vr9Zo0Teumaaq6rivnXGWMKa21pTFm2jTNpCiKkXMunQ/UnFprszAMx51OZyylTIhoMXgzzrvvQSLCo+9mhMXf8zsLl0uLRws2f+5koHHy+ZN/L7rP8d7/rAS6PJ/z9Fd62SDjtHmfx7y56rmcFgycVjF62uuWC7rzu0V+9vrFnSSLvxeFq8WPEMIXRdEURTGbTqfT8Xg8KYpiqrUeB0EwDYJgEgTBNIqicRAEkzAMx1mWTRBxGgRBBQCVlLIOw7BZX19vAMA9e/aMBoPB8UoMBoPzbo77ALe2trAsS7m/v6+jKAqapomIKHbOpd77jIgyRMy01lmSJHGSJOFDHktHSglxHEO73QbnHCAiVFUFzjlwzv2sK6zl/fRtd6W+Kch4W0XeWWOOXCUEOe39b3vfVUOX87ovF+sXWe+bqHB5W+uh25rXVd1WZdRF9++bDK1uYtoPrVLvPOeBi+7/t7WNztqXbuPcdpkWElfZLpf5LjnLVT7z63DTn899P0Zv87v5JrfVff8cLuIy3zerOk+e9Zrl0GPxs+imFgAgCAJotVrQbrchiqKbXmx2PgRHdTu0TEpJZVlCGIarXj7GGHvncAByx3322We0s7Pjsyyz0+kUO50OFEUBxhjvnLPGmMZ7XxHRxDkXCyEi730shIiVUpG1Nh6Px+nLly+TyWQSBUGgvfcKEQURyfmjICIx787nOBRZfsSjb+/F/wEAcN4tznL4cfy/RYCy1F3OawHK8rSWA42TAcpp3tYa5bzvOytsORlYXKS1w3JwsRxanLIsx08uApalO+sXhaXleS9Cj8U0CRG9lNJ770kI4RDRCyFs0zSmKIqyruuCjloHFUKIGSLOELEAgBkRzQCgcM4VVVWVSqlSKVVLKZswDM1sNrPr6+sejlom3fsBzs8yGAwQAOSLFy8CRAyNMQkAJN77bD7OTmatTZ1zkfdezcPDB0sIAWEYQp7nx61A9vf34ccff1ycd0BK+Vo3WIvHxS59WguRs5xWIbb83KJS6azKJUS8cCCxvFynXRRf5qJ3eTrXFZA8xADkMk7bN5Z/v+x2OhEwn3tZLrt/nHdZ3jaNq1bSnnc+1zW9k9O+6bvWH1ql3l1rPXSV/eMyx9xZ87/ufflN0zzP8XvR75KzzmvndZ7vnPMuy5uW7SacXJb78F13HfvuVef7kF3nNj1tm113sH+Zct5Zx/zy86dNd/n8shx6OOeOx+hrmgasta8FImx18KcurwCObmj1ROSXQxAAgFevXkGr1VrdgjLG2DuIA5A7DhFpMBjQ5uamD4LAWmshSRJCRDedTq3WuqmqqpZSzoQQoXMuIKJIKRVYa0PvfViWZfTq1atwMpkEUkrtvVdCCElEx0GIOIKLMGTROgQABJwShMwrHl8LRRARvfeIiDgPF5Zblhy/nn7ewuRn3W2dFk68KRSZT/9C7zltHm8rOL4tDDkRWgAi0vI0T1Tg0Xw5aDn8mI+1QPOQY9HSw+NSU9p5aOIR0RORR0QHAE4IYYmoqaqqqaqqAoBSa10JIQoAKKWUJSJWQogSEaswDCsiapRS9Wg0skEQWO+9/cUvfuHgqND20K++xHA4VMaYgIhiKWUipcySJMm01q0kSVrdbjfNsiwJgiAQRx8MnravPQSICFrr40eAo2OiLMvXLri896dWYrztovJkBfbJC7+T4cdyyHHygvHk+98UppxcztPm/6b3nHzvac+/7aL7PJU+d6my46oVPlepcLjItrpKBfFFpnHZCss3VWhc1Mn97DwVPed13s97lfvodQRJ99FNrPdVA8TTXPT8eHJZzjOtyzpvpftlluWi3yVvOze+bX7nDRLfFBbdhe+fVYUKF3EflvE6zvl3wU3uk9cVgJznvHme4/4iAcji+UX4sfy46LI2DEPQWoMQ4lw9KbCbtwhBlh/n1+wkpTzuCosxxtjt4gDkHhgMBp6I4Msvv6SyLMk55733zhhjtdYNIlZKKWWM0YiopZQaADQiBkSkJ5OJnkwmGhG1EEIBgCYiBQBSKSUBYBGAiHkFr8A5Orrj/TgQWQpAXgs75sGGWPwupTx+HpYCEiI6fh/A62HHchdVZ9UwnxVovKnAd9Z7LnoHz9vCj+XXzO/Kea1lx/L05wWhnwUfMG/psXj/chAyfzwOQuAooHCI6J1zTghhEdF4762UshFC1ADQaK1rRKyklBUR1VLKWilVdzqdpqoqm+e5KYrCOud8EARuf3/f/+///q/f3t5+UGN9nEREuLOzI4bDoY7jOETEuKqqFBFbSql2FEWdKIo6vV6v1e/30yRJAvkOdKgrpQQpJYRhCM45MMZAWZbHF11FUYC1Fk4W3M+qlFk8dzLcOPne5defVnFzMiA5+drTQpLTpnFyud62DqcFNZdx3grHi1aGXXdF5nkqy95WeXCRZbnItC5S6fe2eVxXxdZlwozzrNNlKmxvez1uex4X/c6+quuY7nVt0+tc9+us1D3PtK5zf3/Te962DFf5PC9a4fmm8OE8r7lISHKe4+qyFbeXDX/O6y4HDJfZJy8z/asc2zcdFN6W61yP8+xTl9nvrnKTwJvOgW8qX572PuccAMBx+JFlGbTbbUiS5PjGJbZ683Ojp6MPjpYZYwARqdVq0UcffUS7u7urXlzGGHtncAByf9DTp089ANBXX33lf/zxR6e1tlVVCSGErKpKSCll0zQqCAJljFFaa0lEGhGVlFJJKdW8Gx+NiBIApNZaCiGElPK18EMIIRARrbWCiIRS6jjEsNaKeTc4r/3uvcd5/TAugo3loGQRaiz+XgQeUsqfjc9xVgBy1jgeZ9VLv2ncj9PmgSdabCw771ggp01jqcD6WkCyaO0BcFQ6Wgocjru8mo+78Fr4sShUIaIHADf/sfMWINZ7bxCxcc6ZIAgaAKgRsUmSpCmKwgKACcPQTiYTV1WVOzw89BsbG/7777+np0+f+k8++eQhhx84GAxwZ2cHh8Ohqus6qOs6ttamxpiWtbbTarXybrfbffz4cd7v9/P54OdhGIbqrl2k36QwDKHT6Rz/LqU8DkSKoji1dQbAz0OP0/530nkqjN70+tNCkYu4yHQW63xaJdXbKvtuulLlNl2lQmDZZbbBeUKZy1Z6XnR5z1u5eN5w5rR5ve24Oc+0LjuPk/O5yPyuWvF81rwvsyz32UWD01Usx3n20be99k3/f1Nl5nn2kbP28/Oef857rL1t2d90TJx1Tn3b+e682+A8634dofp9/l67DRc9Xq+z3HCXzpWr2k/Oe1PHTQZ0b5veony9/Lrllh9JkkC73YbNzU3o9/vQ6/UgjmNQiqt2Vg1/GquThBAe5t1gIaJXSnkiokW9AGOMsdvF35L3BP7U/RF+8skn/tmzZ7i1tYXffvstbm5uYp7nOJvNhPdexHEs4jiWxhiBiFIdlYakMUYBgAzDUAKAhKMWIIsusFBKKebBxCL/eO1359xrQcbi9+UWHYvXKaXg5HMnQ5DF/wAAnHN4MsRYDi8ueuP9ogDonLtQkALw5qBDSvnGK4fTmrMuF3IW03bOwfyuEFg0hV0EHQBHH7SUkqy1x78vLFqFCCH84scdbWCHiI6IbNM0VilliMgGQWCcc+Zo8aydzWZuNpu5zc1NN5lM/Pfff0+7u7sEcDTmzAMOPgDm4QcAiJcvX0rnXBAEQWSMSZ1zbSLqeu9zKWWeJElvY2Mjf/z4cbvdbqdBEEillHyXLuwXd5cFQQBKKXDOwWw2g6ZpFvvwW1t+nPz7KhXVJ1938u+TlUDnvcg9a/4n33/a684KQ06b33kr9S5SQXFT++NFK0muEoC87f1nbaPzhmZv278us6438VleZF5vmudl5nueY/C8x9NNuq71vU+uemxdp8ts//OGleeZ1lnzvsh58LyVyZcJnS7yXXbatM5zHrzsZ36ec9Z1ffdcNbS86XLWZbbhdS7TyXLLZVx2ee7aufI6tutVzkuX2eevaxsuny9OK2+ednwSEUgpIcsy6PV68PjxY+j3+5CmKQRBwF1g3RGLEGRxvY5HNyx6POq1gYIguFsHImOMvSM4ALlnliqnT/3iHAwGIs9zXF9fx1arhZPJRDZNI6uqElprGcex8N7LIAiE917OW3CgUkoIIXD5BxHRGINCCLTWCgCAxfOL3+fLhNba10KRk6+11r4WkiyWd/G+xbROWvz/os16l++AOSsEWUz7xPtO3a5vCz6WpvnG/y9CDQAA7z0tz28RiCyeWwQei9cu/18p5efv9/PClfPee2utb5rGdbtdK4SwYRi6IAjsaDSyk8nEt1otNxwO/e7uLm1vb9OTJ09eW6/BYHCe1by3FuFHr9eTYRhKrbUuiiJ2zmXe+3bTNF3vfY6IuVKqmyRJq91uJ+12O1r1sq/CcndYRARVVcF4PAbvPcxDzkuHH6dVeL2pUuis4OG0971pHmdN423vP2v537bsb3PeCrP75Loryq9amXaeaVw28LlqZe5FXvumAO8y77vMtE6+7iLTvo79fJUB9F0IJpddZXtedvmucmzfVGh4U9v6IpWqFzmPX3SdrxIOnWc5bmKa7HxWte0fWpkD4OIhyGWPq5vex992Ew8RgVIKOp0O5HkO/X4fOp0OhGF4o8vFLmYRgCxagCCik1J6IQSFYei999DpdB7egcgYY3ccByAPzHy8EFy0EFlfX6fRaORns5lI09QqpTDLMlGWpajrWmitcT74Oc5bKiAionMOpJRojEEpJdZ1jUmSHM9HCIF1XR+XzOq6xjiOoWkajKLjuuLlFhzYNA0CACz9/zicwDNKlDQfv6Npmgtth4u+fml5LvW+8wqCgBariojknIPFXSBHY5a/3gIlDEMqy/L4EQCgrmsCAPLeU9M0FEURKaW8c4689z7Pc980jS+KwnvvXZIkPo5jP5lM/Lfffku7u7s0GAxoMBi8UwUvOhrzA1++fCm73a5yzumiKCJjTLLo+so513XO5caYrjGm5ZwLvfcPftyP89BaQ7fbBSKCfr9/vL8C/HQH7nnusn/bxeib7q4/K2y5ygXpRSsNbuqO2YdSIXHVyoGbqIi46j7ypule1nWFRKtqlXHR7XnTy/VQjp+z3MT+e13TvO5tf9mg7yy3FTJfZXuet1XKTYReHICsznW2JLguD/1cunCR8sNl3ndVbzpehRAQxzF0u12I4/jCvSSwW+MXNzMiovdHXWZ4gKPr+1UvHGOMvYs4AHmA8KdBspGI4NmzZ35rawt3d3fx008/hVarhXt7e5hlGf7www+Ypil+8MEHAACwv7+PAACbm5vHv0spcTEg8oIQAsMwhPF4fFxCW1TQL4IOAIA8zwEAYDKZHD+3XHEKALAYX+Sk2Wz24K6kjDGQpikBHA1gNxqNjv9eWA5vFr/HcUyL31ut1nGrkOFwCO12m4bDIfX7fXLO0f7+PpVlSdPplIbDIeV57re3t2lra2sRvryLha7FgOei2+2q6XQaxHEcGmMS51zmnOsQUVdKmSNiLwiCjpSyhYgRHHUX987TWkOr1QKlFOR5/loXWOdxlTuF3zaP27ogvcmWDA+l0uE2A5CLuOsVczf5+V/3tO/6tmS3axUtUe7aPK5qlQHNQ/nueZdxAHJ7VnE+Oa3F8aJ1dhiG3O3VHbJo+YE/jQPy2hggi0CkKAqIogi++uqrFS8xY4y9WzgAedjOqvA+Lr3NuwSC3d3d117w2WefAQDAzs7OhUt6u7u7CADw6aefwmQyAQCA3//+92+dzosXL+7+Veo129zcPNeVxscff0yLbr3KsoSnT5/Szs4OAADs7e0BAMC//uu/0rNnzwDgeCwPgHcz7PiZwWCAw+FQzGYz5ZwLnHNxURQJALSttbm1Ntda98Iw7Mdx3O/1er08z1thGEaSb60CgKNu5ZRSEEXRO3uB/K6u90NwHypBGWPvJv5uYex+uEtlCTxlnBB2Nyx3gSWldADgENEvfqSU9MMPP6x6MRlj7J3DAci76fhK66xukOZjQSBcoQJ9cUH37NkzLp2d4cWLF5e2tsPMAAAgAElEQVR63dOnT2l7e/tkwXf5c72OxXsoEABEEASyrmtd13Xkvc+klJ2mafpN0/Sdc704jvNOp5Nvbm7m/X6/k+d5q9PpBFprvrVqCV9wMcYYY4wxxthP5nUfi3E7PQB4770HAC+EcEIIL4Sgpmk49WaMsRXgAIS9yZW+nJcqSflL/ppxwHF+g8EAt7a2xN7enmqaJvDeJ0KIVtM0ORH1lVJriNhPkqSf53n+/vvvd3q9XqvdbidRFEkOQBhjjDHGGGOMncOiO3KPiE4IcdwCxHtPAAB5nh+P78kYY+x2cMUeY+zBGgwGYnNzU/7xj3/URBQGQRAhYuqca3vve1LKtSRJNtbW1jY2NjbWNjY28n6/38rzPG6320EURVJw57qMMcYYY4wxxt5gufsrmI/9gYgOAJw/QotB0D/++GP67LPP+EZRxhi7JdwChDH2IC3CDwDQaZoGiBhZa1NEbHvve9ba9TiOH/d6vc21tbXNfr+/lud5r91up3Eca6UUBx+MMcYYY4wxxs5lHoJ4KaUTQlgAcEIIp5RyzjnvnKO6rinLslUvKmOMvVO4go8x9iB98803GASBBAAtpYyapkmIKEXEtpQyl1KuxXG80ev1Hr3//vuP3nvvvbX19fVukiSRlJLDYcYYY4wxxhhj57LUAsQhopuHIMcDoXvvyVpLAAC//e1vV7y0jDH2buFKPsbYgzMYDAQASO+9juM4nE6nsVIqbZqmHQRBV2vd11pv9Pv99bW1tbU8z7utVquVJEkshBDIo3wzxhhjjDHGGLuARQsQRHRE5ADguAssKaUPw5DH/2CMsRXgFiCMsQeFiHBrawsBQJVlGTRNE0spU+dci4g6aZr21tbW1j788MNH77///sba2lovy7IsiqJQKaU4AGGMMcYYY4wxdkGL8MMLIRYDoFsp5SIEIWMMra+v89gfjDF2y7gFCGPsoUAAgJ2dHQEAstfrqTiOQ2NMKoRoCSE6RJTHcdxfW1vb2Nzc3Gy32xtJknSjKAq52yvGGGOMMcYYY5e1GAR9Pvi5VUpZAHBaa0dEPo5j+u6771a9mIwx9s7hCj/G2H2H29vbIs9z8bd/+7fij3/8o1pbW9OImFRV1fHe5865vjGm3zTNGgCsaa17aZp20zRtx3GczFt9cIs4xhhjjDHGGGMXttz9lRDCCiEMABilVKO1tkop9+rVK5pMJrS1tUXc6QBjjN0eDkAYY/cZbm9viydPnkgAUEVR6CRJgqIoIiFEZq3Nm6ZZs9b2nXNr1tq1uq773vuOECLVWodKKb3qlWCMMcYYY4wxdj8tDYDuhRBOSmkR0SKiEUJYrbX13vuNjQ2vtaadnZ1VLzJjjL1T+I5nxti9RUT4m9/8RqRpqjc2NsIwDBOlVMt73y3Lst80zboxZqNpmkd1XT8yxmxUVdWrqqplrQ2893LV68AYY4wxxhhj7H5bBCBKKSuEMFLKRgjRzFuCWCGEi+PYD4dDevLkCY8Dwhhjt4hbgDDG7iMkItzZ2VHj8VhLKUPnXCSESOu6bhFRyzmXW2vXvPcbUsq1IAj6Sql+u93O4zjOpJQaOARmjDHGGGOMMXZFS11gWSGEWYQg3nsDALZpGg8A9PHHH9OLFy8AADgEYYyxW8KVf4yx+wa3t7fFzs6OqqpK53kexnEcI2LmnOtYa3ve+3Xn3CNr7SNr7WOl1ONOp/Po/fff33j06FGv0+m0wjAMpJR8DmSMMcYYY4wxdlU07/7KSCkbImoAoNFaNwBgpZSu1Wp5AIDPPvuMww/GGLtF3AKEMXavDAYD3NzcFMPhUEkpQ0SMnHNpVVUtIuo653re+773vm+tXQeAtSAI1nq9Xu8v//Iv842NjazdbsdxHAdKKQ5AGGOMMcYYY4xdybwLLKeUMohotNYNIhrvvYnj2IZh6MqypL29PQ4/GGPslnEAwhi7L3D+KGazmYqiKKzrOlFKpdbatlKqK4RYC8NwXUq5TkT9+YDn/W63m6+vr3fW19dbeZ7HSZIESimBiByAMMYYY4wxxhi7quMusJRSDSLWUspaSmnKsrQA4Ou6JgAARHzLpBhjjF0nDkAYY/cBDgYD3NrawtlsprTWejabRQCQElHbe58jYj+O40fdbvdxkiSPELHfNE3XOdfJsqzV7/ezbrebZFkWBkHAg58zxhhjjDHGGLuyxQDoUkqrlFoMft4AQCOEaJIkMX/84x89APjd3V1uAcIYY7eMY2fG2J02H+xcrK+v49dffy3TNA289wkRdaqq6hFRr67rtSiK1vv9/vu/+MUvPuj1eu+FYdgjosR7HyqlwjiOg3a7rYMgUDz2B2OMMcYYY4yx60BEpqqqHw8PD/+/77///usff/zx/43H4+/iOP5zr9fbb5pmrJSqAcA+ffrUISKHIIwxdou4BQhj7K7CL774Qnz++eciCAJZVZV8/Pix2tvbiwEgM8Z0nHM9Y8yatXZNSrkhpdyIouhRu91+lGVZFxFD770UQkillNBaCyEEB7+MMcYYY4wxxq6CvPdERM45VxtjKudcCQCVEKISQtRhGDZlWdrNzU2rlPLffPMNcfdXjDF2+zgAYYzdNTgYDBAABACI9957Tz1//lwDgJ7NZiERpU3TtL33vaZp+tbaNefcehAEa977NSFEP4qiPEmStlJKr3hdGGOMMcYYY4w9POS9d9bapq7roq7radM0s3kIUgdBUDvnTBzHpt1uu++++27R/RW3/mCMsVvG3cAwxu4MIsLt7W0BAOLXv/61BIDg4OAgVkqlANARQvScc2vW2o2maTaMMRvGmPW6rteqqupVVdVpmia21ioi4ltrGGOMMcYYY4xdu3nTDzObzWbD4XB/b29v/+DgYFgUxdR7XwJAo5QySilXFIXf29ujzz77jMMPxhhbAW4BwhhbuXlYgV9++aX453/+Z/n48WPx5z//OYjjODTGxHVdJwCQWWvbiNgJw7AXx/Gac27DGNO31uZBEORBELQRMYajcxsHIIwxxhhjjDHGrh0RkbXWNE0zPTw8PJhMJvtlWQ6ttVPvfYmIDRHZyWTi/umf/slvbW0Rj/3BGGOrwQEIY2yVcDAY4M7ODn700UcCAOTjx4/VbDZTQoiwruukKIpUStmy1ra997nWuheGYT+Kog2l1DoA9JqmaUkp2+12uxWGYSSllMidqzLGGGOMMcYYuxlERNYYU85ms/F4PD6s63ospSyUUpWUsiEiq5RyAOCBu75ijLGV4QCEMbYquL29LTY3N0WWZeLFixeyLEs9nU6Duq4D730MABkRtcuy7HjvuwDQj+N4rd1urz969Ohxq9VaD8Ow2zRNhIhRGIZRnudhFEUcgDDGGGOMMcYYuxFEBEIIJ6VstNYzrfXUOTfTWhdCiDoIgmY2m9kgCBwAcOsPxhhbIQ5AGGOrgNvb2+LJkydyNpvJFy9eKCLSzrnQex967+O6rlPnXBsAOkSUI2JPa70ex/F6u91eX1tbe9zv99fiOG475xQRSSmlDMNQBkEgheAhjhhjjDHGGGOMXRvy3oP3npxzzhhjnHMVIs6klFOl1EwpVUopa621ybLMbmxseA4/GGNstTgAYYzdJhwMBggAotfryW63q6bTaeC9D6SUQdM0SV3XKRGl1tqWMabrnOtGUdSLoqjf6XQ21tbW1vr9/lqe52udTidPkiQFOB5HBBARuPEHY4wxxhhjjLHr5L0H55yrqspVVVWVZVnOZrOZtXYKANN5S5BCKVWHYWgQ0ZVlyeEHY4ytGAcgjLFbMRgMxNbWFg6HQxEEgUzTVJVlGSJi5L2PvPcJEbUQsWWMaRtjOtba3FrbjaKolyRJf3Nzc2N9fT3P87ybZVmmtQ4QUQAAhx6MMcYYY4wxxm6M956qqnIHBwfVcDicFUUxNsaMjTETRJwqpQpErJVSTdM0zhhDxhgOQBhjbMU4AGGM3ah5ywz88ssvxd7ensjzXDZNo621gXMuJqIEAFIiypxzHWtt1xjT9d53iagnpexGUdRrtVq9fr+/vra21u52u6nWOlBKyVWvH2OMMcYYY4yxh4+IqGkaOxwO6+fPn8/G4/GEiCZZlk3CMJwhYqm1rojItFota4zxk8lk1YvNGGPvPA5AGGM3YTHGB37++eeY5zkOh0OVpqlyzmlrbYiIUV3XibU2a5qmBQDtpmnypmm6xph8EXzEcdzt9/vdXq/X7Xa7eZZlaZIkIQAIHuicMcYYY4wxxthtICKy1vqyLJvRaFQMh8MCAGZCiJlSahYEQem9b9I0NVVVOecc7e3tcQsQxhhbMQ5AGGPXZtHa49mzZwIAxIcffiiklDLLMqmU0pPJJCKiiIjisixT732raZq29769aPkx/+mkadrpdDr5o0ePuhsbG61+v99qt9tpFEWBEILPXYwxxhhjjDHGbpsHAOO9r621hRBi6pybAsBMSlkgYlUUhTHGuLIs/aoXljHGGAcgjLGrQSKCZ8+eIQDAzs4ODodD8eGHH0oppex0OkJKqaSUWikVaa2Tsiwz730KAC3nXAcAOt77LgDkiNhFxDYiZmEYtlutVve9997rPHr0KOl0OnEURZq7vWKMMcYYY4wxdtsQkYQQXkpptNa1UqoCgBIRCwAoiKiUUtbee6u1dnt7e7S7u8stQBhjbMW4+xjG2NsgAMBgMDg+X3zzzTf45MkTfP78OX7yySeQ5zm+fPkSrbVibW1NlGWpjDEqDEMVx7FGxMA5lxhjWtbaVtM0HWNM23vfFUJ0gyDIwzDsEVHHOZc2TZN0Op10c3Oz9dFHH2W9Xi9qtVqBlBIXVrc5GGOMMcYYY4y9a4wx5vDwcPynP/3ph+++++75/v7+d865P3Q6nd+12+0XcRwfIuJsfX29aJqm/uqrr8y///u/W0TkEIQxxlaIW4Awxk5zHHp89tlnsLOzg+vr6/j73/8e8zzHX//61/i73/1ObG5uorVWTCYTDMNQKKVEWZayKAqdJIn23uuyLANEjIgos9Z2vPcda23XWtsBgDwMw7zb7fZ6vV5Pa90GgNhaGyRJEnW73bjVakVxHGutNbf8YIwxxhhjjDG2KiSldPMWIJVSqgSAUkpZeu8rRKyttaYoCleWpc/znLvAYoyxO4ADEMbYsuPgY2trCwEAPv/8c/EXf/EX4rvvvsM8zzGOY4zjWHzwwQfSGCOstcI5J6y1UgghjTFKCBEYYwIACIUQgXMuQcSWMSYnonwegHQRsReGYS/P895f/MVf9FutVqaUCr33QkqpgiBQSZIorbVY6VZhjDHGGGOMMfZOQ0RCRC+lNFLKSkpZElFBRKVSqhJC1EmSGKWU3dvb89vb28StPxhjbPU4AGHs3XXcjdRgMMBFt1abm5uY5znOZjOxtrYmAEBMp1OZpqmM41h47+XLly8lAEjnnPLeK0SUQghljNHWWu29D5qmiYgogqMQJInjuJPneS8Igh4AdJ1zbSLqdDqd9traWjfP826r1YqDINBEhIiIQgiUUqIQgru8YowxxhhjjDF2q4jIE5Ezxti6rouyLMfW2hEijpRSYyKaAkAJALVzzgCA6XQ6bn193QMAhx+MMXYHcADC2MPzs7CA6Kdy12LA8m+++Qa3t7dhd3cXNzc3cWtrC7Msw+l0KjqdjsiyTHrvJQCoNE2lMUYTkTLGKOecJiINAJqIAmutJiJNRIH3PvDeh8aYmIgi732ktU6zLOt0Op1+t9vtaa073vuUiJI4jtNer5dmWZbEcRxyV1eMMcYYY4wxxu4C772fd2s1m81m48lksl9V1YH3fiSlnAghZmEYVlLKJssy4713o9HIP3361HPrD8YYuxs4AGHs6s7bOuG6Cj+nzm8RciwCjoXFGB6Lvz/99FP8/e9/j5ubmwAA+OGHH4o0TbGqKhGGocjzXDjnpJRSKaUUImoppUbEoK7rQEoZSClD731Y13VERKH3PnDORQAQAkDonIustbH3PjbGxACQImK30+n0Hz9+3Gu32xkAhESklVI6DEMdRZGWUnJLD8YYY4wxxhhjdwIRuaZp6sPDw9HBwcGrw8PDl1VV7TVNs6+UOiSiWZIklTHGKKVsHMfum2++8f/wD//A4QdjjN0RHIAwdg5EhABH4cLW1haur68jAMDTp0/hq6++wm+//fbUivuPPvrouNDz1Vdfwccff3ypQtBiPou/T5vf//zP/yDAUcABALC39/+zdzc/chzn/cCfeuuXednlUiIlxvYvjpD4QAO5CDCQQyDpGCRX+phj/Gdo9W/4TxCvuRmIpVMAJ0QOgXlQHEGOZK24szvv/Vr11PM7cHo9Gs3uzpJLcil9P8BgXrq7qrpnt3uqnq6qkSIi+vd//3fa39/XRERJkqj5fK5+8pOfqKZpdFmWSmutiUhnWWaISE8mE0tExlrrYoyOiJIQQqq1TmOMadu2qYikq8BG6r3PYoxpjDETkSxJkrzf7+dKqR4R5cycWmt7b7zxxt7+/v6tW7du7Q8Gg5611sYYjdZaaa2NMUYrpRAAAQAAAAAAgBtBRCIz+7qul8vlcjybzUYickJEE2vtXClV5HneGGP8/v4+f/XVV/Hx48dCGP4KAODGQGMjwAVWgY+zx+PHj/Xx8bFO01QlSaKcc2o8Hisiovl8rt544w06PT09235vb0+IiG7fvi3ffPMNERG98cYbV/4h5JxTRERdXuv5vfnmmzSdTtVisVDWWmWtVUVRKCIia61q21YbY1QIQRtjlPdeJ0lyNnl5XdeGiEwIwSZJYpqmcVprS0QJESUxxlRE0hBCtgpypCGEjJnzGGMWY0yZOfXeZ865PM/z3sHBQX84HPastTkzO611OhwO+2+99dbgzp07/V6vlxhjMNQVAAAAAAAA3Fje+2K5XE6Pjo4+/9Of/vTHo6Oj/3POfZOm6bG19jjLspExZsTMyy+++KI9Ojriw8NDBEAAAG4QBEAAtlMiQg8fPtR37txRd+/e1b1eT8/nc5OmqT46OjLWWpUkiTbGqNPTUz0YDM42Xi6XlOe5EBH1ej1ZLBbEzNLr9YSIiJkv/TG0v7/fpaX29/dpuVyqboiosizPXneThNd1rQaDgZrNZjqEoLXWKoSgrbWambW1Vtd1bYwxOoRg27Y1RGRExHjvnVLKrub5cDHGhIgSEel6e2Ra6zSEkIUQUhHJmDlj5mw1/FXqvU/7/X5++/bt3v/7f/9vePfu3f5gMMiY2SilTJIkrtfrJXmeJ0mSGKWUvu4vDQAAAAAAAOC6eO+XVVWdPHny5LOvv/76f4+Ojj43xjzp9XrHSZKcaq3HaZpOQgjVaDTyDx48wNwfAAA3DIbAAvgudXh4qFbzZhgi0iEE84c//MEqpWye56ZpGlNVlXHOaWutNsbo2Wym0jQlERFjDMlqUo7RaCRJkoiIiPdeiIhijJf+IDo9PaU8z8l7r8bjsWrbVmVZRlprJSIqxqjatlWrIaQUM+vZbKZWAQ6jlNJa67MeHl3Ag5kNM1sRsatnR0SubdtEa+201mme51mSJHk37BUzp6vJzZMQQjfnR7oKhrgQQhJCcL1eLzs4OMhv3749ODg46O/t7aVERCKitdbaWquttZoQfAUAAAAAAICbKa6w974MISxjjHOl1Mw5N1NKzYwxc+fc0jlXn56ehh/96Ef86aefCoIfAAA3DwIgABsODw8VEWki0nmeW+ecmc/nNsborLVuPp87pZRlZhtCMCJirLU6hHDWqG+tlaqqxForMcaz19576QIj1tpLfxgtFgullFIhBKWUUmVZKvU0sqGaplGrOTOU914bYzQza++90VprZjarQIhhZhtjtMxs6WmvDycijpkdETlmPhvqKsuyrN/v94bD4cA5l4lIysxn6zOzW6WVdK9DCDbGaLMsS4bDYba3t9fb29vL+v1+8oK+JgAAAAAAAIBrJyIxxuibpqnrup6XZTkNIUyJaGqMmVlr51mWLbTWhda6bpomfP7553E19BUAANwwCIAArBER9fDhQ/XNN9+YPM9NVVWOiFyMMVFKpW3bpkVRpN0E4UopS6veFSKim6YhY4wQEWmtRWsdY4wiIhJCiFprWfUQkaZpiIjO1l/HzGqVhgohKK21WiciZx9477WIaGbWImKY2WitzWroKcvMtgtUrMprVz04XNezg4hSZk6NMZlzrr+/v7/31ltv3cqyLDfGuBijEREtIjrGaIhId5/FGM8e1lrjnHPD4dA55zDHBwAAAAAAALxWmJmbpqnn8/l4Pp9/M5/Pv27b9jiEcEqrIEiSJAtrbZllWfPOO++Ed999NxLm/QAAuJEQAAH4M/Xw4UNNRObWrVs2hODSNE1FJG2aJieiPISQe++zqqpSpVSyCh4YpZTpghKrwIc8jVM8pZSKq89it5yZzzLWWp/9UIoxKiIipZSKMSpjDK16gehtARCttXbOmSRJbJ7nxjlniciKiIkxdgGPswetBUC6Ya26QIgxJhsOh/3BYLDX7/cPer1eZq213WTwIqI2X6/Ko/68K1qvhgbDMFcAAAAAAABw461uXIwhhNi2bV2W5XI+n08mk8losVgcE9EpM8+cc0ulVFlVVX3v3r2GiPzf/u3fMoa+AgC4uRAAAVgREfr1r3+tDw4OzHA4dFVVpYPBoNe2bc9732fmgfd+wMw9Zs5o1WtiNayUXQtIkFJKlFLS9fjQWkelVOyCIusBD2b+VgBkNazVtwIgRKRijHr1sRIRpbXu5tLQ/X7f5nnuBoNBkqapc85ZETEiYkII3WsbY+xeu9VrF0JIYowuhJBordPBYJAPBoNhnud7WZZl1lr05AAAAAAAAIDvLRGJ3nsuy7Ity7JcLpfz+Xx+OpvNTubz+ShJkom1di4ihbW2unXrVk1E7f3794NSKr7q8gMAwPkQAAFY+eijj9QvfvELTUTOe58OBoNeWZZ73vs9Zt5r2/aW934/xjgIIfSYOffeZ0TUza2hVxOSUxf8UEqJMeasN0j3TETU3SHSrd+Vo+tNoZSi9V4WXeCjm/dj7bVO07TrvdHb399P0jR1IqJX62lmPhvCSimlu9erXiLdHCFGKWWdc241CbrTWqMXBwAAAAAAAHyvhRBiWZbtkydPlrPZbFoUxWnbtqfMfOKcG2ut58aYgohqa227WCwYw14BALweEAABWLl//7768ssvTZZlLs/zNEmSXCk1UErti8iBiLwhIm8Q0S3n3CBJkl6WZflqKKmzIbCMMWc9OlZBkLMeIV2gY7N77GrZt8qzNtwUrQU/aH3YqS4Ykud50uv1ev1+f9Dr9dIsy1y33WpILdWlSavgybZnWg1hZYwx1lqjNgsFAAAAAAAA8D0TY+S6rtvJZLIYjUaT2Wx24pwbpWl6miTJWCk1E5FiOBxWTdP4Xq/HDx8+lF/+8pcIgAAA3HAIgACsPH78WN25c0crpcxqSKiUiHIi6scY95j5QCn1ptb6jTzP95IkGWite6seFN8KgBD9OfjRvV5/7qwHQrbFGtbm1jgbGmstWHEWDNnb20sGg0GWZdkgTdM0SRJ3vUcHAAAAAAAA4PspxighBF8URTGfz+cnJyfTvb29iVJqkqbpTGu9zLKsDCG0g8HA/9///R8/ePAAQ18BALwGEAAB2DAYDCiE0M25YUTEikjCzJm1tt/v94d37969tbe3t59lWX81pNRZL4r1QMZ6wOPplB3nd49dLd9qPRCy3hOEnmZIaZrawWDg8jx3xpjzEwIAAAAAAACAb1FKRWutT5Kkcs4tnXNzpdTcGDNfzf1RNk3T3L5920+nU75z507EgAkAAK8HBEAA1ty5c+fstdZahRA0Mxt6GghJtNZZmqa9g4OD4d27d/cGg8FAKfU0srEWpCDa3qNj9fnWIMhFP542017/TClFxhjlnNNJkhhjDH6FAQAAAAAAAFxA/izGGFsRqY0xhbV2kabpzDk3U0rNY4xLrXWZpmktIj5JEh6NRkKY/wMA4LWAAAjAFs45iU8J0dNgQ4xRa62tcy7p9/vZ3t5e79atW30ieuU9LrrgCe5AAQAAAAAAALhcjDEys2+axtd1vazreh5jnBljptbaqbV26pybaa0XvV6vmM/nzWeffRaIiI+OjhD8AAB4TSAAArCmrms5ODiIIhJFhI0xgYh8jDEQESulIj29y0NprVXn1ZYaAAAAAAAAAK6CmbmqqnqxWMwXi8Xpcrk8bprmRCk1zvN84pybhRCWRFQopWrnXHtwcBCIKP7qV79CAAQA4DXxyu9cB7gp7t+/L3/9138dnXORiNhaG6y1rVLKxxi9iHhmDiLCMUb23scQwtNuIiLo/goAAAAAAABwg3VDXjFzDCG0ZVkWp6enk5OTk9HJyclxXdcnSqlxlmXTNE3neZ4vq6qq8jxvZrOZf/z4cfjlL3/Z3RgJAACvAfQAAVjTNI0YY1hEAjN7EWmIqFZKVTHGhpmbuq6bxWJR93q9WmudZllmkyQx1lqNziAAAAAAAAAAN9Nq2Cv23nNRFOVisZjP5/PT2Wx2UhTFyFp76pwbJ0ky11oX3vv6rbfeaj7//HMmIj48PIyveh8AAOBq0AMEYOXx48cyGo3i3bt3w97eXisiTYyxJKKCiJZKqUUIYVGW5fzo6Gj+xRdfLL788stiOp02TdPwqhcIAAAAAAAAANxAzMxFUbTj8Xh5cnIyPTk5OV0ul6O2bY9jjMcxxhMRmVhrZ0qpcm9vr/nqq6+YiPjBgwcIfgAAvIbMqy4AwE3x29/+lkajkaqqSoUQVFmWioh0CMEys/PeZ8yctW2bLJdLV5alCSHYPM9Nnuc2TVOjtUZQEQAAAAAAAOBmECKiGCOJiNR13S6Xy3I0Gs1PT08n0+n0uG3bJyGEY6XUyFo7stZOiGgmIsV0Oq0fP37sR6ORfPDBB7jpEQDgNYQhsABWlFIiIvHRo0d8enoaiKhl5ibGWMUYC6XUgplnIYS+9z6tqipJki8fBk0AACAASURBVCQtyzJh5gwdQAAAAAAAAABultV8H+y958ViUcxms/lsNpssl8vTsixPiOjUGHOqtR4rpWbW2nmapkVVVU1RFIGI4uHhISr8AACvKQRAAL5NPv/88zgYDEKapno2mzVKqTLGmBlj5sw8izHm3vtEa52GEHpE1CciJkyCBgAAAAAAAHBjxBgphMBlWTbz+bxeLBbT2Ww2LYritGmakYiMlFInMcZJkiRTY8xcRIo8z6sQQtu2La+CH6jvAwC8phAAAVjT9QL59a9/HYuiCD/+8Y+bqqqcMaaIMS6cc9MYYxpCSKy1mbV2aK3dN8awUgo/iAAAAAAAAABuDvHe83w+r4+OjmbT6fS0LMtxjPGEiI6TJBlprU9jjBOl1CzLsgUzl4vFopnNZv7o6Ag3OwIAvOYwXwHABqWUHB0dcb/fD5PJxBNRba0t8jyfaa0nxphT59zYOTfWWk9CCNOiKBZFUZR1XTfMHDAhOgAAAAAAAMArJ8wcvPdVURSzxWJxWpblExH5Wil15Jx7kiTJSZqmkyRJFsaYcm9vr57NZp6I+MMPP0TdHgDgNYdJ0AG2+OSTT+if//mfKc9zqutaiYiy1iqttY4xKqWUsdbaPM+TLMsSa60jIqOUUtZaq7XWSin1qvcDAAAAAAAA4IdKRMR7XxdFMR+Px6dFUTzx3h+nafpNlmXHWZaNlFJTa+08SZLlrVu3yqqq2n/8x3/0P//5zwUjPQAAvP4QAAE4x8cff0yPHz+mEAINh0PK81y01qSUIqWUcc4ZpZRlZts0jQkhGK21TdM0cc4ZrTV6WAEAAAAAAAC8OpGZy7Ztp/P5fMTMR0qpo1UAZJTn+amIzI0xS+99Za1t/v7v/z4QUUTwAwDg+wFzgACco5sP5NGjR3x0dOSVUrUxxoYQLBFlMcY0xpiXZZkwsyUilaap9Ho9RUQxTdPUWmuMMZow3BwAAAAAAADACydPcYwxeO/rtm1nIYSpMWZsjJl0Q1r3+/1JlmWzwWBQjcfjJk3T9quvvmJC8AMA4HsFARCAC6yCIPzo0SMiIjo6OjLD4dAsl8uEiGxd166ua922LRERW2tZay1N04S9vb1Br9frEVFiDDpbAQAAAAAAALxoIiLM7Nu2LcqynFZVdVxV1TfMfKyUGiVJcjocDsfW2tnt27eXy+WyNcb4qqo8ETGCHwAA3y8IgABcTj7//PM4GAw4yzLftm1NREWM0VprnfdeKaVi27bh9PQ01HXNBwcH3nvPWmtrjLEGERAAAAAAAACAlyGGEJqiKKanp6dfL5fLo+Vy+XVd10cxxhMimhHRkogqpVRz9+5dPxwO+YsvvuDf/e53QkQIgAAAfI8gAAJwCaWUHB4eyr1792Ke5yHLstZaWzKzISJjjBFmjnVdx6ZpYlmWxMxirVV5njutNYlIZowxq8nRMRwWAAAAAAAAwHMQEYkxSgghMnOMMUatdRSRpmmaWVmWo/l8/vV0Ov26aZpvmHmktZ5Ya+fMXFpr6zzPfVVVfHp6yqPRSA4PDxH8AAD4nkEABGAHh4eH8vHHH8dvvvkmvP3220pENDMrYwwppSIRcdu2XNf16jeXpizLdJZlViklMcaY53nmnHMIgAAAAAAAAAA8nxijtG0by7L0TdP4EEKrtfZKqapt2/FisTiezWZH0+n0G+/9E631Sa/XmyilFsxcDQaD5q233vJEFP/jP/5DHjx4EAm9PwAAvncQAAHYjTx48CA+fPgwfPPNN/SXf/mXipmlLMuYJElQSvkYY3DOxRCCqutaTk5OpGkaLsuyffPNN/2bb755WymlkyTB/x0AAAAAAADAcwghSFVV4fj4uBqPx0VRFEvnXOGcWxDRiff+qKqqr4no2Dk3staOtdYzY8xiMBhUxpiWiAIRyS9/+UsiBD8AAL6X0BALsKPVhOjx4cOHwTlHTdPIm2++KUTEVVVxjFGYWYmIjTHScrmUuq6jUoqMMarX69lVjxFljNFKKQyHBQAAAAAAAPAMRCQysy+KohyPx/PJZDIxxszSNJ0450YxxuPVxOcnzDwlopnWehlCqKuqar/66iv+m7/5m/iq9wMAAF4sBEAArkApJUTEH3/8Mf385z+XqqriZDLhXq93FgBRSpmmaYSZJYQQnXM6TVM9GAycUkoRkcqyLDXGYDgsAAAAAAAAgGcTQwihbdtyuVzOxuPxiVLqNEmSkzRNR9baE2PMKM/ziXNuJiJLpVR5+/btumma8P777/Or3gEAAHjxzKsuAMDr6OOPP6ZPPvmEDg4OxBgjeZ5LVVWyCpCIUioqpUQpJWmaKqWUijFSCIGUUtpa68xTCEICAAAAAAAAXBEze+99tVwux2VZntR1/SRJkidpmn6T5/kTY8yJc26cZdmMiIper1cyc3Pr1q3wm9/8Jn7wwQcY8goA4AcAja8Az2AV6IiHh4fy3nvvCRHJYrGgXq8nzjmp65rruuYYIxMRVVUVnzx5wiGEVikVkyQRpVQQEY4xaiLSWuuzobG01uqV7iAAAAAAAADADSBPRWaOIhJFJCqlYgihEJGZMWbsnBslSfLEWnuUpumTJElOnXMzpdQiTdMiz/NqOp02X3/9tX/06BEfHh5i6CsAgB8IBEAAnp0cHh6KiMjDhw/l9u3b4r0XZqbhcChERCEEijGqsixjjJGNMSFJEur1eiQivm3blpmdUspZa22WZc45Z7XW6J0FAAAAAAAAP3giEkMIoWmaNoTgmdlba1tmXnjvp0R0bK09TpLk2Fo76vf7oyRJpjHGpYgUzrl6Op229+7dQ/ADAOAHCAEQgOfUTY7+ySef8HK5DEVRtNZaQ0+HmFMioqy1zMw+hNAsFovWGFPN5/MDpdR+27b9NE3zPM97t2/f7u/t7eWr7QEAAAAAAAB+0JiZ67puxuPxoizLZdM0S+fcUms9Yebxcrl80rbtE631E2vtCTPPrLWLEELV7/ebvb09f/fu3fD73/8+Hh4eYtgrAIAfGARAAK5BFwR59OhRePTokUqSRMUYKU1TYWaJMXqlVNO2bbNYLFrvfUVEixjjrRDCfpZl+/v7+945p5IkMdZao56OhbWaN50wJBYAAAAAAAD8IIiIEFEUkdi2bVOWZTkejyfT6XRSluXEOTe21p4S0bhpmtO2bcfOuROt9dQ5NyeiIk3TpixL//bbb4evvvoqPnjwIBIRAiAAAD8wCIAAXBOlVPz444/V0dFRuHfvHiVJInVdx8FgwMaYRkSqEELVtm09m80qZi6YeRljLAeDQR1C8L1ej5xziogoTVNnrbXOOf2q9w0AAAAAAADgZRERDiF4731TFMVysVjMJpPJaPU4McaMnHMja+1YKTU3xsyUUjNjzEJrXbRt29y6dcuPRiP+6quv4qeffho/+OCDV71bAADwCmCYHYBr9PHHH9NoNKKf//znUhSFaK2jcy5679k550MI3R0nopQ6m7zNGCNKKRIRxcyKmZUxRltrddcb5FXvGwAAAAAAAMDLwMxtVVXlfD6fzGazk8lkMprP50/atj1m5pEx5lgpNdJaj7XWU2PMTGu9IKJKROqTkxN/dHTEeZ7H//zP/5TV0Ffo/QEA8AOEHiAA16gbCouIZLFYSFVV0RjDZVl6731DRGytjTFG6SZFZ2YmIm6ahsfjcQwhSNu20RgjqyGxtNZaE5HGcFgAAAAAAADwPbEa6Yokxnj2WiklbdvWVVXNJpPJ8Xg8PpnP5ydN05wy8zhN01Ol1KkxZmytnTFz0ev1irquq4ODg6aqKt/v98Mf//hH+dWvftUFPRD8AAD4gUIABOCaKaWEnv6Qk4cPH8o777wTkyThL7/80u/v70cRkaZpiJlZRIL3PohIG0JovfdeRJiI/HA4DHmes7U2JkmSGGMSrbVBZxAAAAAAAAD4PogxxhACt23LzByIKGitQ9u287IsR4vF4mixWDxZLpcnIjI2xky01lMRmVprp0mSLKy1FRE1/X6/uXv3rr9//37o6uWvePcAAOAGQAAE4AVZ7w3y8OHDWFUVExENBgNSSsXVkFi1tbYSkYKIliGEgpmrpmmK6XRaaq1LZq6Hw+F+nufDJElSwtB1AAAAAAAA8JqLMZL3npfLZTObzeq2bYsYY+WcK4loXFXVcVVVR977ERGdGGPGSql5kiRzZi5CCEWWZZUxpu33+22SJOH+/fuslIqvet8AAODmQAAE4AVa6w2iPvroI7l37157cHAgSin23vsYY22MqY0xpYgUxphaa90wczWbzaq2beu2bYNSSowx1hijtdbdXSyKniaulFLUDY+FYbIAAAAAAADgBjkb3mr9WURi0zTtYrEoj4+PF4vFYsrMsyzLplrrUxE5bprmWCl16pw7NcZMnHOLGGNhjGmUUo0xxnvvQ9M0/Hd/93e8qoMDAACcQQAE4CXoAiGHh4f0s5/9TKqqYq01hxBCr9cLIQSvlPKr+UBCjLEty7L13rfWWu73+9E5F2OMe1rrhIh0jNGIiBYRrZQySZJo55xZBUkQAAEAAAAAAIBXTkSImTmEENq2ZSIKIhKVUr4oinq5XC5mT5167ydJkoyttWNr7YiITolo4pybpmk6JaIiTdOKiAIRhc8++4wPDg7iP/zDP0QEPwAAYBsEQABeosPDw9jNDTIYDMhaKzFG6fV6IiIxhCCrMVB9VVUtM7dFUYT5fN4qpaokSfaVUlkIIRURx8yOmZMkSZJ+v5/s7e2laZqqp3OmAwAAAAAAALxaMUbx3oeiKKqiKKq2bRsiapRSTdM0xWKxWNR1PW3bdlzX9XQ10fmEiMbW2qm1dp4kydw5txwOh9VisWiGwyF//vnn8ejoqJvoHMEPAADYCgEQgJdsdVdK/O1vf8tPnjxRt2/fVtPpVKVpSkopEpGotfZa61YpVZdlWZ+cnCwXi8VEa73PzANm7jNzL4SQM3M+HA77d+7c6TnntLVWO+cwTwgAAAAAAAC8cquhrvxkMilGo9FsuVzOmbl0zi1jjMu6rhdN08xjjFPn3MwYM9Naz40xU2vtwjlXEFFBRPXR0ZEfDAbh3Xffje+++66shoBG8AMAAM6FAAjAqyGffvppfO+998IXX3xBMUay1kZjTNcduDHGNMxchRCqxWKxKIpiIiJ7Mca9EMJejHHAzP0QQp+Z95IkGQ4Gg6C17hFRZq21Wmuj0R0EAAAAAAAAXrC4EkIIvKK1jszsi6IoFovFeDqdjmez2YyZ58aYOREtRWQhIgtr7VwptdBaL40xS631kpnLXq9XWWubPM/b4XDo//Vf/zW+//77giGvAABgF5gnAODVUYeHh+q9997TVVWZk5MTm2WZHQwGSVVVqYjkIYReCGEQYxyIyJCZhzHGPSLajzEOmXkYQhju7+/v3759e+/tt9/e39/fH+7v7w8Hg0GeJElijHGvekcBAAAAAADg+42ZQ9u2frlc1lVV1d77VmvtRaRummYxGo0mo9FoPJ/Pp8w801rPtNaLVS+PpYgskyQpRKTUWtda6ypJkto519Z17e/du+ffffddVkrFV72vAADw+sAwOQCv0CeffEJ/9Vd/Rfv7+3Lv3j0uy5KNMdy2bej3+14p5a21bZqmrda6TZKkdc611lpvjPFaa6+UCsaYQEShaZrAzFEppZMkcc45a4xBTy8AAAAAAAB4oUIIoSzL9vT0dPHkyZPJkydPJovFYrxYLE4Wi8WoLMtjZh6JyEmapifW2pMsy06zLBtnWTZO03SaJMkshLBUShVEVKVp2oQQ2n6/H37zm9/EDz74AL0+AADgStADBOBmUCJCH3300VmPkOVy6Xq9nlNKpcycW2tz730vxjhQSg1DCIO2bfeYecjMt7TWe9bavVu3bh3cuXPnzttvv/3mYDAYZFnWExFNREYppa21BkNjAQAAAAAAwLOIMUZmjszMMcYoIpGIove+Loqi+PrrryfHx8fj+Xw+d84VWutCKTUnopmIzJl5obVeaK3nWuvCGFMMBoOCiOq2bdskSVoiCkQUusnOHzx4EDHfBwAAPAvcGQ5wM6xP3hZFhD/55BMmojCfz0O/3/cxxiZJkpqISu99ISL9NE3n3vshEc2993ve+z3n3DLP82o+n9cxxr2yLAfMnCilUmtt2uv1sjzPEwRAAAAAAAAA4KqYOdZ17YuiqNu2bZm5Ncb4EEJZVdViPp+P5/P56Ww2m1prF6vH3Fq7TJJk2QVFtNZLrXU1GAyq4XBYxxjb09PT8OMf/zj827/9W/yXf/kXXs3zgaAHAAA8MwRAAG4gpRQdHh7G9957LzjnhJljWZacpqm31tbe+8o5t4wx5jHGOTPPkyQZxhj3RGRRVdVyPB4vZ7PZvtZ66L3vO+cG/X5/+Oabb+4754xzDnODAAAAAAAAwJUwMxdFUR8fHy+Xy+WyqqrCOVcS0TLGOK+qaiIikyRJptbaudZ67pxbKKUKESmZuRKRWilVhxCaxWLRxhj9T3/60/D555/H//qv/+KjoyNB8AMAAK4DhsACuLnU4eGhun//vqKn8/WcPW7fvm2LokiVUmmMMWfm/mqy9KHWei9JkgPn3IGI7IvInvd+mGXZ/nA43P/Rj350cHBwsNfv93MRUfR0+K2zZxHR3XuttTLGaGOM0VorteqmAgAAAAAAAK8nEZEYo4QQeDWUlSiluoADrQce1j4/e18URT2ZTJZ/+tOfZpPJZFGW5SJJkoVSaqmUmjPzrG3bKRHNiGjunFsQ0ZKezulRiUijlGqbpvFpmnqtNRtjOM9zfv/99yM9HSEBgQ8AALgWaMwEeA0cHh7q+/fvq8lkog8ODhQRmTRNbb/fT4qiSImoR0Q9Zu6v5gTZZ+a99Uee5/u3bt269eMf//jg4OBgv9fr9URExxiNiJju9eq9VkoZY4zNsszleZ4kSYJ5QwAAAAAAAF5zzBy991yWZVPXta/rmpVSUSklWuu4CnpEpVRcvf/Wo6qq6vT0dPnVV1/NTk9P58vlcu6cWxhjFtbahTFm4Zybreb5WBhjiizLlkTUEFGT57mn1Rwfo9EoPn78OBJR/PDDDxH4AACAa4cACMBrQkTURx99pO7fv6/u3LmjNidKb9s2E5E8hNAjooGI9Jl54L0fMPMgTdNBmqbD27dvD3u93tBam4uIY+Ykxpgws4sxOmZORMQRUdrr9fLbt2/37t692x8MBom1FsPmAQAAAAAAvMbatg1FUTTffPPN8uTkpJzNZrVSKmitWWvNSik2xgSt9ebDr+b6qJfLZTkej4uyLJdN0xTOuaW1tjDGFMaYwlq7NMaU1toyTdPSOVeFEPzJyUl45513/HQ6jXme82g0ksePH8vh4SGGuwIAgBcCjZkAr4m1O2Hk8PBQERH94he/IGOMJEki1tpYVRWnaepFpBWRqq7rMk3TRdM0/Rhjz3vfm0wm/bIse1rrjJkzZk6ZORORNMaYhhCyGGOqtc739vb6xph2OBxGY0yWpqldDY9Fq+GyFK0FUrtlq/KSUkpba5V+ighBVwAAAIAbYW0InBhjFBG5tobHa0wKfgB+iHf87/o/ctmx2VzevReRc5cRkTRN48uyrKfT6Xw0Gi1Go1GllPJdkGP13FprvdbaE5F3zjVa61Zr3YpIHUKomqapiajSWlda68JaWxljKmttlSRJFUKo8zyviahZDXsVvPf83//933xwcBB/97vfIfABAAAvHBojAV5f6uOPP9bvvPOObtvWxhitiNjxeJyISKKUSr33aQghVUrl3vsshJARUUZEWQghJ6JMRHIRyZk5V0plIYRcRHKlVP/g4GDw9ttv7/3kJz/Z39vby51zbjVElloNmaW7OUPWAyNERMYYba3VeZ67NE2Nc04TzjkAAAAAN0IIIYYQuCiK4L1n7328pqTRkAlX8joHQM4LZFy2T5vbXbC+bFu+/r6bn6MLemzO49G911rH1XrStm07n8/rP/7xj7Mvv/xycXJyUhBRq5Tyq0BIa4xpjDHt6vPWWlsTUWOtrZVSDRE1SqmzBxHVvV6vNsY0RNQmSdIMBoM2TdP29u3b/vj4+FvDXSHwAQAALwsaIwFeYyKiHj58qN955x19fHysl8ulJiLjnLPWWtu2rWNmR0RJ92DmVGudikhGRDkz5yLSizHmSqmcmXsxxh4R9Xu9Xn9/f39w69atYZZluTEmYWYbY+weZhV46YIhZ5OoJ0lier2ee/PNN/P9/f10NVQXzjkAAAAAN0DTNGG5XPrj4+NysVi0ZVmG60j3OnuSXOZZGs7RO+VmuWnBj4vKs7ls299SjPHS9ZVS3/k3Weu58Z1Ax3pvjvVnETmbuFwpdTZxuIhIF+zo5u9YPZ8NbxVC8HVdN6PRqDg9PS0Xi0W16t1xFvzQWjer55aIGmNMrZRqtNaN1rqJMTarkQfaGGMrIm2e594Y44mInXO+G1LLGMNffvllPDg4iA8ePIg37XsHAIDvNwyBBfAaW/1wjIeHh/Lhhx/yw4cP1Z07d9RoNNJpmqokSUyM0dy+fduWZemUUtYY083zka6CHlkIoRdjzEQk9973Yow9Zu5rrXtVVfVijD1jTCYiaQghjTG61fwhTkTOgiGr4IcWEZ1lmdvf30/SNB1kWZYnSZJsBEDODYasD6W1tq/Xcsw2035VP76vq9v7i87/RZfjZeeJRo8X60XEOLedD26K5ynbq4wHP+8xRSz7++lVX5d28Szn8FdZ3ufJ+2Vcr9q29WVZNqenp8uTk5NmNpv5Z03roobe5yzmlfK9zHrjNDx1Xd/Rs/7Nvoi/kef5ns8rzyXl/NayGON56599th7o6AIcG9utP5/Xq2M92BFXQZCzScuJ6OxzrXUwxgRjTFBKBRHxzNyWZdlNSt5Ya88CINbaxlrbGGNarXVDRK0xprHWNs65JoTQKqXaEIJv29aHEIK11hMR53keT05OYr/fj5PJRFZBj67c3zleAAAALxpqsADfY2tzdJgvvvjC5HluiqKwIQQnIknTNGlZlpmIZDHG1HuftW2be+9zZu4xc87Mmfc+DyFkzJzGGNMYY0JEaYzRxRiTLggiImb10L1eLzk4OEh/+tOf9u/evdu7detWop7ektSdd7bOH7KaK4RijJuBigvPV9363fY7HJfnrXBdedv1/HapmGmtz83jorvLdnDlsq+XZZeyP+8dmddZGb5q2a/Tq2h4e9UBg/X/wc3/42e16z5dtWH+WY7VNe/fM2+/XvZdznubnqfsu+b3Cv4WX7vftbvcTXzdeZznea9Lu6T7sq+7RNvLvOu14Krlfd7r2HVdr3bNuygKPx6Pm//93/9dPnnypBmPx+Eq21+UZ1f+F3kdvEra38cbIK6zp80ux/KydZ73N9Z1/q287ADItmDG5rZdmUT+PN3O5uebvUC6IMf6Yz3w0d0Mp7WOIsLda/pz4IOVUlFEuJvbg4jCarJzvwqIeK21d861xhhvrfXGmNZa26Zp2qz1CPFa66bf77dpmp4NlWWM8Xt7ezyfz/n+/fu8KiMijQAAcKOgBwjA99ha9+p4enpK+/v7MpvNZDAYxDzPeTqd8mqM1zrGmIQQuqGyUmbOutfdwxiTKKUSa23CzKkxJiGirkeJ7QIh6unk5y7G6MqyzKbTado0jVNKdfOAqKfFUyrGqLTWZ8Gap7/l1WbD2beCJUTfCmKcvd9slNvWwLe+XlfJWK8kXaVxZ1vFc73Cc9HYvtsqR7SlcWetInRu+tsqZBeVY1vZtdZyUWXxecp+WXrnlfOifb1KnX9bo8yzNOKtb7+r58nnWV2lYftZGs7Py2czras0fq8HLrZtt/n/flE6u+Z7WZrb0tkM0F6U12WBkouCulc5tpcdu408d1rvsnW3Ff2i723XvK6yzTnpvHYBEKLLg+O7NApedE68bPvzzqvnnOt3Pg+fdx06r6G8c9F5c9t197KgwWZ+3fqbDfTn7c+ujbJrv7ku/ax7fdGyrozPch3Ztk/b9qOua57P5yGE0GitQ5ZlvLn+8waLrrOR/qJ8dnEdRXmVPYq2ucrx3fV33lXXuerfyrPkcVXP+11fNQiy3nNjW/BvPdDRnRe6bda37YIam8tWQYyz4a2659X3H40xZwEQWusJQkRRRNgYw10QRERYKRVWAQwWkdA9YoxdcCQopQIze611YOZgrQ0iEhaLRSCiYIwJzrlwfHzMv//97+OdO3fi/fv3u0ANAADAjYIACMD3nFJKDg8P5f79+/HOnTvy/vvvxy+++CI655iI2Hvf5nluyrK01lpb17UVERdjTFY9PJxSyimlkm74rNXrRCmVMHNirXUi4rogCBEZY4wVEbtcLl2M0RpjrFJKi4heNVJ1z12vkLOAiHr6q349EHLW2LjeANm97tbtXq/t+05DbnXH6ZxF32lY2Vj3O3d4XbTtZkPNZYGEteVbK1HraV5wl+22YMNF+V4YzNhskDmvPN2669tepWHronR2aRQ67+7TqzQoXUfDzcsOgjxvr4RdAxkX9bpaC2ruXMb1/+fz1t2W1y49IdbT2DyPXLTdZlk2zzPr557NbS4LyG5rrF/P77z93tZLbtfjfd4x3nRRQOKy72A9z6se113KdoGdglHPE2C5qosayjZd1Ih/UYPgLj0GdjnnXdCAee714LL96Na97Hp13vXjnED5udeJ9bQ2rzvbro+bAZ7zjtNlPRnWt9nl5oL147ctv6vcoHBR8Gzb38Zmft57qaoqeu/ZGBOzLJPL0r2oDBfty2bezPzdDXb0rNfVm9RAf12uIwBy0T5d5e//ecq2S1l28azn+F3/ji9bl84Z4mpbMOS8nh/rgY91q3PB2esu+KE2hrpi5rPPuvda6y4Awl1AZBXk6HqHcAiBkyRhIuL4FFtrOcbITdPEJEnYGMNVVcUsy7goipjnOX/22WdycHAQP/30U/nggw8QAAEAgBvptbxTDgCeiTo8PFQffvgh0apHxePHNahYxAAADKNJREFUj/Xx8bFO01T1+31dVZWpqkozsymKwhKRaZrGGmMsMzutte2CIs65JMboiChZBT+cUsrGGC0RmRij1VprY4whIqOe9v7oAiCaiDStgh6rgIfuGvFEpGutOguGbPQUOWvwW2vY+tYd2ZvrXtYofF4FbrPSsyVo8Z3KzbZG//UK5GZjz3ojwOa662XbvLtslwaezX1Yb3DZzOeyIMNFd7ZtOw7nrbutAWwz/Yvy3dyndRc1sKwvY+aXEgS56T1ANm1rlL8sj6f/4n92UWP8+nYXpbFt3YvW2basK8tmWuvnjcuCJ5vH0hhzaTBl8/N1lwVfzguArO/ftmDGLg38m+fB8wI167bt/3nrXFCGc/+mzivDszRgXXSev2kBEKLzG6SvEvzYvJ50zguKXNSAub7elobpC4MS29ZbX/eyYP955+lt15Jt18N15wXdtzXEb8t313TXnXeN7pZ1+ewaHOrKtv5+87fCtvzP26f1z7ddk5i5G5LnSvt9XhnWbUvzon25btedz8u+pp+X33nf83l2OQ67BKjOy+u8bZ/leD3PMb6GG0AuPN4X7X8IgYiIjDFnr7elu758PV0RkRDC2ev1z0XkW4GP9ddt24pSKiZJEkMIUSl19gghxBijdO+999E5x0mScNM0MU1TZmap6zpqrWOe52yMid57eeONN6L3XtI0jXt7e/Lll19KlmWxKAp566235O7du3GxWMhoNJLHjx/L4eEhAh8AAHCjIQAC8AMjaz0qiEh98sknajgcqjzPVZIkajQa6cVioUejken3+zrPcx1jNFVV2bZtbZZlhpldjNGlaWqVUrZtW6eUssxsich0D73CzGYV+FDds1JKaa31eq+PVeOr2ixnFwBZb5xdbX/2mujbFZ/NdS87LrtW3rdVgjYbVi5bZ33ZZgXzgkDGpXlsazDZLPdmWa5SrvX327Y7r4J40R27F+XzLHeO7pL2VSvmzxMAuUo+1+F5K/+7/K/s0ih+XjrnlW8zjV0DJdvSu2yd9bJdJQjTrbMtz/UAzWXfwS7npsuCH5tlOW+dzay7F5cFfs4ry3ku+rt5nn28qvPyuskBEKKLz1ubyzc/f55G8XU7NJDuEgS5sLH7omvDLmW86Nq1bluAe9u1cZfr6Hn5n5f25j6dd01ez3+Xcl20v8YYISLabHTdlua2cmymtS2di3T5bxNj/M6yZ8njeVxnXhft64tw3ne1uU+7lGuX47CezlWO27ZyXrT9yzqOzHzh+X6Xcqyv472/cPm243fZ+cR7f7Zd978RY5TusxijWGslxigxRmnblrr3zCwxRsmyLDKzaK3PAh7dc1EUXYBEtNaxC3ZoraMxJrZtK8aY2DSNGGNiWZayt7cnBwcH0gU7lsulEBFNJhP52c9+JqPRSFYTmhMRJjUHAIDXAwIgAD9gXUPQRx99pD788EN6+PChevDgAf3617/WBwcHqigK3e/31f7+vmZmE2M0ImJijEZrbUXk7Nl73/X80MaYs4f3/uwzZlZaa0V0FsDQXWDDWktKKdVVVtaDGsysugbGzQa/yxozL7tDfNNmZWizAretYWKzMr/eULGtcnVZw9R6WusNG5uVrPPuMDuvAWf97rRd93fbet0dauvLrbVyXsXwoor6+jbW2u+Uq1t+USV110r2eXldZlsDzlW8zAaTyyr7l+n+Py8SQvjOOs65ncpj7e4jb65v273ezGfXsqynZa39TrmYWV1Wtu5cct56m3mcZ9t+XbTNtoDA+nlvc7vz/gbWt9m1rOflv+m8wNCmbWVbz/95/n63fa/XncdV7XLeepZz8La0djnPXNTwfVkAZP08eF5e5zXSX3a9uqhs266H28pw1cbWbY2TF13HzsvjsuvyZcdtl+/7siC8MWZruTfT2eUa2H3etu1FWV5Zl+555XzRrmN/rvK74Trskt+uZdp1/5/1+98sx2Xbv4xjue33wbOWxTknTdNcuHyXNDfTWD8/dGk0TUMxRuneM7M456Sua0qSROq6JuecVFVFzCxJkogxJiZJIswsIYSzR9ebI89zadtW2rYVa22s61rKshRjTDw4OJDFYiHj8Vju3bsnjx49or/4i78QIqLVfB70+PHjs3J++OGHCHgAAMBrCQEQANhGHR4eqt///vfq5z//ufqnf/ondXx8rJfLpd7f39f9fl+PRiMzHA5N27Y6SRJdFIUJIWjnnGZm3ev1FDNrrfXZcwjhrBeH1lp1nznnaNUZRBF9u9LCzKp775w7W5YkybcK3KWz/n49jfMaaIkub2Q/ryLjvf/OsvXKzC6Vqsvy7pavp7Ut3a6yuW3ZeY0e1lo5r5K6+flmupuVPaLzAwVXCSCsp9s0zdZ8tjmvYrqZ3rPYtQzfF977K/82SNN0p/QuWm/Xsqyn8axlXd9u/VyxeV65rCzrQgjqou3X81jPc/31ReepzXXX09tlvS7tXRuF1l0WNLis3Jflu779dQQodh3K7VXadv24yGZQeJvnaVS8rGF68xp12bXmsjJ1dzHvWqb1htmLttt2Tbto/c3z+7Nexy661lx0DbmOa9eu16jz1kuSRIiI6rreJZlzt7/M895M8DyqqrrW9NI0vRG/C3Y99lfd/13XPy//y7Z/GcevaZqdrgO7lCVNUymK4vkLtdLNtdMJIcj6sqIoKMsyyfNclssl5Xku8/mciIh6vZ4QEc3nc+r1euK9l8FgIJPJhAaDgXjvpWma7n9aqqr6Tm+Od955Rx49ekQHBwexC24cHh4SXTIfIAAAwOvsxlcQAeDV6oaievjwobpz544aDofq+PhY53mulsulTpJEJUmiqqrSzjllrVVFUai2bbVzTg0GAzLGqKqqFBFRXdfdXdSq1+sR0dNKSnfn+fpnXRk2KzFt2yoiojzPv1PeXe5gvw7bKvLM/EyVhfMqX2VZXrh8XVfZvGzdi5Z3+V1mM41n3e9NeZ6fpdNV+HbZbrlcXkf2l5bph6L7X30RBoPBlbfZVp71dK6jvN15iYio3+9fuO4ujSrdeWwXuzbSnLfutvPgeXq93pXyuyzv67S+H905/nm8rGvBs7hKQ/B6A+N1N+Luatt1Y/OzXa8fRLtfry4rw7Pmf156z3ot27x2XbR83XVcu65yjeoaTs/TNbBet36/L7PZ7IWk/bL1+/3v1W+C6XT6XNsPBoNvHY/JZPJM270oy+XywuvAyyrHpr29vbN8T09Pv/V+NBoREdH+/r4QEb3xxhtydHT0nTSqqpI7d+7I5mfdcFVET4esIiI6OjqSrjfHgwcP5KOPPiIiIszbAQAAPyQ3tnIIADeOOjw8VERE9+/fV0REd+7cUUREn332mXr33Xfp888/V4PBQBERPXnyRP30pz8lIqKf/vSndHR0dHa+OT09/c65ZzKZqLfeeus7mc5ms53PU2mavrRz2t7ennSVlOfVVXLO8+TJk53TOjg4eCkVmTfeeOOF5HPv3j0hIvriiy9eRPLP5Mc//vEPpnL41VdfvRa/C7pzy/p55WXYdu56mSaTyTPlv+3celVXORe/anfu3KH5fH5jy3ud14+X4bJr1LqbeL06z3Vex17lteu6rlH/8z//cx3JwGvkD3/4w3Nt//bbb/9gfh9dp3feeefsuD169GjrOj/72c++dWw//fTTby3vAhrr1oMbnVWQYx2+MwAA+EG6sZVDALjxng4AuzE09UcfffSd88qHH374nY0fPnyI889ram3iwxdmswIHsG7bOeVlwbkL4PX3oq5juHbBD8mHH36IxvSX4AqjOuL7AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAACA/98eHBIAAAAACPr/2hcmAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAIBfE7oLmOab5rgAAAAASUVORK5CYII="></image></svg><style>@media (prefers-color-scheme: light) { :root { filter: none; } }
@media (prefers-color-scheme: dark) { :root { filter: none; } }
</style></svg>
